��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�V=�?�"n;-܃��E����g�Q�\��c{��aO��x˖���\�� =���{��H7
v�����ǂ�n���P�{�q�h�m�h()���On�xA�ͧ[�Q/�L��5o#���/+�>��{9�rp���<z�ɠ+Yz��a�X�Ϸ4G~e�vM��]����9aQ9�"��W���N׳�NUzo/���mD��2���2q�Iާ��0��p=k��	)-����:�ݫ�-���QT�uG,�%��b��N0΢N�
�~D�t�m� �T���^���}�s	��W-����F�΢W�=�ވ��L=��+eKr�:����H!=�G2�����u��� %�(�Y9���-7�XW�t�'����Q2d4��()�7�H/۪<��<u��΁��2BPl�#��4U}D�'<���'��?�7��y�i滖(�J��]lp�+�x��ZY��B�,�xP@��]�oן7��"{��<�Գ�Yh�3��-:����@.T�tt�&�IG&�rށY��8Qw�IYz���?��؃m�rܯ��,[� ���W���r�ħ�� �l"�Ke�͞l�@Q�f���+��h�TV�P�5֤yq&F���.��K�C*}�Cҹ���`��U����
�%gb�.V�=�ŀ��ꁺ�U����ݿ���C���hWI�Y@��Q1 �-4Xەm��\^$u�,"d���u��+d��j*w�Ŕ>_&��Q!�ae��U� ��߱��2$!&OQ�f�E&|+�M�~�/S�&
e�ȼ;��
Ʊ��F��y��W?��_[w��S���Ƕ��û1�S��Z�{~��5ɦ ��~(�Z5��,I�ු��k�ƶQ��Kw�0�v������,�q���}�������sP��Kw]��jG����8p���a�奏��D4��:l������}��T'(BSh�x��;���F�#�j�$��(�կ�t4ȭ�8�� �..2jZ��٦U�`��m"@�t�)X>��N�H<u�t�oH�����∟�[A(K �B��ť�������΂��&�S+��1�=��`�}7���4Mg�f	*�7ѧ~���U��̇�
8O�/�@�G��J�����v���|4P�A	=>�^G�(d�v-�`�|�-"V�yo��C?/�����/^tѓP	���O��ޭ�3���]0�Q�f�y��
��)R�9�$��ΰa�B
h�n�~� �df"��,�xS��{).]t��0L�,�-�֗w���M~Lh��"��`�A��C�����[vu(���z����P@1<��ӵ���u�C��y�޴��)�Q�[�[�jnf0�c�`nyB�)��]-)g��~YR錽�B����tI��:�$���mo\a�uL������._wzT��Ť7���1pA�+�"�ږ�uTm���B�#���ECѤ+`�5�����<H��O��OQS�ڽ{��_����q8ɀ�$Ꞧ|y��c��_L��k�w��p>I�J���)�hd��W�~��#\3�[.b����fU���*y���<禧��RAm�I	̩�/0E�9/����l������L�5��k�:<'����!�-M,�ܽ�	�<|���Y\*���g|���Q!1g8�/�=����9����$�>��i�lk��l�m`݊������uP��'���L�{�H�:���2l{���e�(�8��0��pC�Y�9�z�����B*��y�����oQ�F߄�D���v[.5^ж|{=2�m(r�7!k+�q���a��9��e]80���XY���@����<�{�xb�Pd�_)*��P��E��:k�;$�䦭k��mθ�����=b�qo]H�]��et�]el��$
�vZ��+KS��~mQ�Ǿ�!���T�
g �/R�:�[ވm@���#=�c��]���n'4wC��`7�?a̍������4���q���~��L��V̇~vڍ�iNԝA�ҧ���w�#��#�%��1Ցbm^��׽����su�ب�hY򭡽���!�D�s�C���uK�Z�sչ����X��GE��X)YBa�'hF�sN����|;Aĩr���땴���
�"����Ў���iTF/\v��r�ݤP@YA����D����/4�M�D�'�R��F�q���p�W��\��=�����Ä��ι��Հ�lb��0��3� �>�^��V���ic�U�\c�~És��0`�)�\�d �2��۫�A���-H~�K�ÞB:�қ�h���N��W`B��1_պ��``��'y��s��.�)j���RA�:�∜���"�p���:@� �8L�)y�&|�dK^.i!��b0���J��e�qmt4��w�D�;���ʥx|ӧS-��t��[>�����4�Q��ϳ6R��A�ٲ����At�t1���2�m���k��!5�
�)�·�w�.}�I/�Қ�xƎ��'��sH��.�D]���~��R�������2���7�CpPɄ	��T,�K��kۂ'F����&vN�a�W�e�`�Q����P�=� ��,\���,F�X���	V]�i
_ϴ&�5*�ˠ�����jY��٭�\�=�$Ɣ���*�f���%�fbT~P�H)��yw~ܽm h��L�iP�P��*���wi��p���:��۝Iٲ<�"����N����{�dG.^�	�qI5��l f�` �+s�A��ZO��9��@�N%{�F^�[�gQR��8�N�6���j�Rb�/^Vn%G��^���m\�A�l���OW��9�����0�7sz��,<�b@Y.���$v���m�ݡ.ǒY�Ϡ����a$�H�z|���d���,��zp���4��B&��r����_	/�c#p9�]>�&�v���a��Ǐ�)+`e�s0�`϶�Y�/hm������ H,0��<�w/���C~=+��P���S/�n;e�؄�]��g�Bk�S^wӡ�(Z�f|g��̕�q�������������}l.�H6�2]�oFJ�Bc\L�Q�v�C�k��J��Þ6qC�n�C��Bt��Ѻ*Vܛ��U����ԮS4��4�n��J�P��L��P�Q��s4k�;�M�n ��+A�~Xy5,�9o���2���`kqP�1�/9��V=z]������o��9Oj������7Qh��s@U�ʤZ\�ڤ�N�<�!9��t��M��>E���"�=b����X
t��('��7�I, ����5e4�A8���L=��v�
��[&�	Ϸ֜��+�Cl��hn1�Z�w��-��1Z���%�$�-��[>�ˑ�8U��%�Ԫ �~���\�y⻬ٹ��l�d x^&��Z�om[[���E(m#D>�����c]q�_�. ��*�?��
A�{"�,�g��w��t~����@��#�s�1�YF�WJ	�m��x�3��Ȱ��Tk�g��;ͯjTt ݕ̦ ���H���&%�/�j��Q�I�^�d u�k�
<�����Ӫ�����N���z�Lg��զk�SѶ���^���аgrsO�F.W�FO�΢޴���r��Z6ӎ�- I�Ϻj*V��
On�V�pB�[/���_��]qYH��m^�ҹ��N��8{�bi4y���u\���t���e�y�+����������t��S�d�� ��)�~���gy����5�x������$V}~��1؜4T(B���ˁ�gP��ܔ�Gq)�^uiSA��O�@��e�(D6���J ��e�"�}����U�Hh�Ǚ��ch�P[>����I�Z`�fܦ��2�,�z�͘��o�S��)VdAp��kg�So���E��h��C����0����L`���U�/�g#�Z��k��8 7�ZR[1G��Ц �O+z���fo�M^����{I��C�.dM���Y� ��f!/���Y���A>�D���ǐܪ��%l�R����SրaK���v@.�C+��)���| ��ZE��g��5{�ƀ�W��˗A��AHG��Φ�%� nL�)����N{�z#\7�A~s}��2�1>d%�ҥV$%���ɔ���;}lή���M�j���a� <\d��S�ɇ��06+)���e���w ���������ey��Luc�+��r�eX�K׫�􄋟�c��,�1�=�\##���3�Aq���'�6�AX}�)�:Z|�eum�?(r����x��q���~�h��S^��ŵ"�t��Hz��$��H`nn����Ϯ�e�9e���W���)���$�*4ìT�C���d����⻺�$�R�a?3#�BjQv��\z�~ �H"���1z�ף&����o)��(oX^��so�V~�n���B���Z��n��ˀȧoa��Gȇ�Z�(+MإA����b�Dl���Ń�5��Sݯv�W�%��;�,���*0���[�{�|���YAR����>?�l�% R.��;p��yHڙ=�"[��d ���X�X:�����k�x����.&�1�W��o�ƍ�]c+�>{4վA�������P:L� �|D�.c���n	���	Va(y��|M֮�q���v��2� �WgH�����Yz��~p������/q���8V�'�Őg��I��1h���-���������`Z7Ga0c������K�5eIҝ�_J}��Y=j���E�����!╆�����~b%�:si�
�n�7�+���6hFO����5����)
�5�՗>�����~���'<��蔇7 ���*K���D7W_������1
 ��
���S4j_���F��ţY�Q��@ʭ6i>Jq�� 3v�)����\W���G��P+fW,ŶZ[�����y� p��	J� ��fͲ��V�mH�1����f�F�0�!1�*���Nx~c�#�����_��~tiVSh{�3D��40�	����IYG}�7'J�T��H�ߩEl����@�,�g�?m~��_wV���n]:�{�q��f�7�eh�l�z�ΫI��b\أ�F*%k��/j:����Iҙ�6 %��PBSfn���@����W�4�پ����u���&�'싩�J��W��:G�⬢V�U�`�ŵ��H�=7P4J��Ӏxsd�U��Ø���:�"4���n�2��֩�8����'��)D�p4�}�@��Y��\�K���-����eӢtQ�~�Y��ڬ8�B�u�����]5�����9�#�����������]"����gC ����|�Ǡ/j�B"��8`U	�6��2��!&!v�ց��߷�����R���w�S��9S����"s�4M�R>�|XN��w8��2�#ʲ��J1e�N�_qe��׫3�l��X�l����b2;%汸����@X9�ku��۷�� ���]�KHp���'v���+"1��=���)�n�c�J^��nYVh����N�Yը��[T��*��x�ִ�3�'�U��&91��>�^�s �G�¢0���+P��4���-Zn�o�H�3	(��D��GZ}td����Y�O��P�����g7t�j4\N���*�$�9M�"��HR�)��E�7tlF
|�%�3�?��"�y��ʫ*�T%��w�a��\k�)0���� Ɋށ���㄂����R�2��� }%&� ��mF$���� �̽��S}>��߿��;y�@g�ԩah���92�
>=]�܅����F!�&8����3���x1Gz���4��ֆ��N2r�e�e�qgs1�5`���డ�� �d�ӸZrL��@�3Ya�|�RɈH�q���}�͊gI���}D/�̨�ζD˹��n_�QB?-��	��Չ�zǰ������만{@p��y�(��m��E
I&�[·��j�vq��d��r��OΚF1�t�������#7�e�=@âv,�z1�Qw* ��2� �u��ot��LA���������9���MQT[�zGd�����A��J�Bf����c$GЂB?�\Nƒ�0�c���lQ��~� ǴXel|:�l�e�.o�� �O���81��E�^Cm"���)�>�;q6-�C�~S������;մr/֭��!]�+R#�|��;�9z��WM	{���e��^�}����9�2��k��#*o�!|nG%�o��(�mq@�{�xOY��|6���D��\]���Kjw�H�lH+<D�]��iB����`ִ��G=��r�f�B��f�4�n�ٹ����W{�����O+ %K������e�Z^+u���h�}��=��ؓ��n+�*����bAz�-� �n��z�4n�b��MhJ#�_ck�������O%X	�������u��x�7��W(�r@�6��}��N�z�r�e��q�$>�=�?�')c,A��y<,nqL�%�s�ڂ�������j�#�_�͚�e^�:�=e��u�D���G����[Q���eA���-����R�4�V�bc�fЛ�PL?�5	�ƨ�g񫮺mXN���/l�������56=
�L��6�'�\�׶��J[@W��d�i�܈���tn�@�J�`����.�߇���:��-���˰R]z4�<��{�ׇ��	oG!��q@�O�8�d-�F��,Փj�y�6}_�Fʒ�(fC��C!�Z�	>��-���F�B|+�z8^�b]֬h����)���F ��ؘp�/-�?>(�^r�4���;U�:�}Uń�(Z�T�fk=YEE���5�*o�	��Y����(MXo���ط�*���&�9�jH�)����l,6
y�~�@��o�bQj��
�h|���I��3cՏ��w��k5 �
v�>��t�:{�+]�}u;���g-�QF0���i�v=<Yj|#j�]��%�-8l���昡��gj%J�OP���Ѯl�� T�ϩ-����S��炗z��#ƅF�[�5
��E�����ŏ(z��COp��]�l\�|zG1�)�8�MQ��1�<�	|ްd���
�L�g/a�%���0�)θ)7D��+D�g���j�AE�`��c��)���J�r�&�� �n�8̽��uq�㔗��UA�=�d���*nN�{[j1.����ZV)�ū���ߣn��E� �#e0��M`>=5��4��J�h��_{0��\J >u���a��D�"/���y�LE��[�o���T_xj������[։Գ��u��
<�BS�Qh�T���Z��g"��I�������Er��pms*�tײյ<;�o��_�O61Ý����{G�	��R���#)(B�&����p�k�nh����\�P��-8�C4Q�/�H?EW���V4�S�0�$wd�psT�&HH}�h���&���CZ��34�t�qACPĀ	�7��=G?C�x�����A�*�޳H�|H��y���y�n,쿯_
���I�/j�j{�2>J���Ҁ�0�K	E������ >W �	H�I0-F��dެ��@9�6�z5:����9���1��hB��-���Ab�3MG�	��l
��a_�����<0L�y���m��vo���R��ӆ���"���dh!(w�*Πc��W@��&Wc����SZ˷{	d�~s�P����!� ��>5ԇ�d���qm�l��S�����F���t>\B�v�*s��D��a�ch���vc�g��v�.��kH���M��AAC���� 0�'�T{`Q��t2ރ����2�.�'+ܪ	D1U�M*uI�zat[9|Gw�@&�3"�Q��s�')sër�y����U�xA=8>$=�	:�c��&�Г�Z�gg(����S�� �i,��w���81�c����q@���孪o�Su�y��h�T���_�P�u2���+�I��=}�����0+�97U�J0�y��XYA[#;|���i���S�N�?����R�\���<�T����g4����m	ر�aK$�5��Sݒ��S������8O��	�6��8	��I�W��ӵ�_��3#/D���u�g�K����'<oA�;�ߤU��ʞ�����0�L��B}��{������E�����v���Up{���Y׭cp� q|��Չ��F"�b��߼?�3tG1�u'�5~7_"	���yzR:�v{~�Z�s��؋	��QC����^^�M{X`h,���-T��۱���^��O2�������2~�wQ���.q�&�����g�)L��K@��,�o�aވ�yM�ަwg��#rK_��.�a]h	�>Y�()/��=�f$���|p�?w�>#r�r"��9�|󹔱�X�C��|Xԣf����ś�{iOKP�&��lU׽��f{��s�/�D�<��,c�ƩcZ�˘�9T���������V띜0�qe���t�Qb�#z��zi.⢢�_�\��k��f� ��$)e��z��*Ͻ��F���WR��X�0[RPMI�e}�w3��%��ɠ!�"G� ��uŉ�����Sjtڥ]K��Ƶ�Q#�7F���d{��.�ى��)��%U�� ����T�J���D�O&8��
Nּ����0��7�S�[Zr ��k�z9���jUd@Jn�zKHZ~ӭ
5�̀��<W�F'��}Aw��I_��z�>r�&d��`	>�����C�@��o�����84���6:ks�v�V��2˽8�_{lʮUr�&�]v���T;N�θ�-3D~^��������zZc����T�5F�����3�E�ٕ��Бs��a�3��~�����4�p�"��2���O)�oMȿ��o�kwK.��<(X��l��8����j������}�j֜�t)�
���P�;���h���,�R����3���?���"��g˜�s��X���a�b�j����ϱ߻G�S��L:�#Jia�u�G�����9
�������H�5��Q��.�H�CyE�\��Yqe�
��Hd��Q.b�����1G`��l�*��̼��
O��=~���?�"ie�w�xV�����@�n���l�	4Y��;�O�\i�l������)��nW�����WK�VNV�lI����/İTB���<`�vt��B�ɚ,]922}ܴ��N#F�D����.��6�&��<`�.�E�&�-5���i�q�J Lƭ�{QZ��'�?�����?n@(7���q��j�Zy�sǨw��&[^����޲�����/�9��LĶXч�*�m� ���S>�����UӇ����=i��� |�|-�މb������{�d�2�$�J\�DiǨ�D��l&���
l#�>ŗ���es�YOŖ?W��.���v�kZϷ��Ɂ�`��1���ы+榥RϷ�μR��"I<�%t8�׽���>�/���W���AT��6#J��,�1�(W���o�y�����ز:(��q'�(K�]!��z�v��{�.N�����(#��S+:@Z�򽵱Ä�4���[U�b��I�
�$&-�K�~0ӝ���t���@Y�Q��-E{��c�j�A���P�9�>�-�����L�o�g�I�4(�G�x�*%�P"�]�s��D�BH��i5o�S�g��\(�^�@ܐ]�mQ?$���b�:�
����Z�:� ~�wx&�F�Q��e"��M�S��6#� H�#u1݌m��e�ϕ�Xjƿڨ����_)~6��0��?��Ҿ�Ƀ'L�,���ݎ���9X�`�pq�/���4��Y&)_��	5� ]C#�����U]�{XP�m�)�wO�L8����5��3�)�:�!B�Iy	l�fLg�"�T��~�=�x��f��Է�����YsghWx����e�`!*�ƏJF,����+� ���Kn�^� ��Y�G�ҼM"/����JzM3��J��Cww�J����ؙ�8	�*L�n��9��e��Ď;p#<��� ��r�S|���R	�vѳE�õ�d,J��=�KY����'��,�q>+S*!C��u��AzAZ��׳�����b�Ց�[�a����qc�bb� ��vy��V��+ ��
�w�1HG�Ƌ�Hq�RC�N�v��y%����*�������6N�g�s�Z�5��di�:�u�8m�����V��w	�֞DF��g��a�'��0UCd��'�lSGM  꺃�����y�m�@9]c$1�C��R����n��� ִ�����d�o��ȷ^ _ �u'
�]����5E�{ʌއ��ĝ*c4l5���j�E����G�Y̅ͨ,����\2�%�C�nÕ]h˼���!�(!ʂ�{��x��Cr�~��$>���
���aU	�`����v�y	
���'�.,|(��Ru̟�TFs`��*e�e�{���b�D�����h�Ď���U��*�e���D��)�
�O�mo!kI~�*�i�ǡ���ګ�:,�@�W9�@Ƞ*[�||n,�X1�">�_���RMD���]y`�,�Mͽ} �h�Zfo�H�|&
�v�&�������"|G.���Zt�B�M��y4�df�!�����
�6��U��&�*�����2C�a/{H��^�/D`��ՠV��F�����z�	�FN�bVNr�ac�Ą�p�/F�A��TKB9笜F��ͩ̎y
]�Β�_5zR�ó�?]�Az�d
ƌ�z�q#�2��7� �bLix�4`�)�β��fnL��<���ͭ�r)H�T���Mov�wWS5���X#^��(�b��R�}Z$[E.���S�1��H�k�*�3'	Jh�E�,KS2�^�xfiu�����t1 F4�&~� 8�(8�Ϥ�#�m�?�g�Qd�[���!��F�����oFW��&��9�����֧����d߶��Q�GKz�yWV4�6�*X�E�R�@#��H8�ء�U�IƂy������1���ͩ���)��̮l���/�`^LQ�9�K�aL�.|狽�k=�i��n� ������&�Ȣ�,z�~eڴ�D��P�1/��F�ndA�V�m�zg�|L�5ud�!��]bvj;H�Xa�<�j�ya7.R�B�( �*��Z�iOPp͎��
��6�-�bJ����^;_pK�*nx�s�\��b@�����	�B��|�~k�"��GR!�|i�Q3Ud��{��&���D.�*������z�/M������N���I޶���R�W���O_��J�i�SkK}��E�y��XF[;.X��I��)����z 	�GG���p���2����Y@��DyV�_�	�6P=��S��ۭ�]�ř6��a	�%D=�wR�I��Fѿ�p��&�zMբ?���^d!��t �t�C���Tz�ߠ��q��jN�EWU�	:+;�8���{��K��N���*�'�T����f�,y4�@f�VO���c�P�K��u�:D1�M�~���=3�|].�����@WThM����
������V-�$�:%E�o��?����(�TY���Y_�G�8�|�%�e�c��Ь>��0>�{���g��*ցx��T��㣀�&��Sb��'v����) �Z�䱉Io�[ӈ��[K7'�}�k��oשVa��\����]��p��soʄ�J��)UQ�K�����?�j���s7�􁎂b���_A����pa����ve���3]�/�����`��`�,��� ���G�pͽ]�su���{���p�.���c�qλЧ��8�����/1G�Y7�`�Y�GR�J�pJ�����6�O)1�ޏ�:�1�,�u�EpLidu}i�u�o�	�.c��#�)[a�"����i� �_V+���=�׶��j��-�ͻ2.�
�|�A�v�!�����d�޳�,��|52�H�wD�-�5S>�R���뉼˰��`��p��`��1���G������қK�Q�.`.2����Z�l�آ*a�}���B|T�_!FeS����̎��_-\u\l��x�B�^������	��Ūe�#<���Cq/��⟕��YZ�"(ɡ�]i ������'�Y���%U�����.�V&C�k�&]�vl/�v���Ԛ��fr����`J��Z꟩�O����oܱw�6@5���&��̵��d3�1n�\��hm�@뼸���*�ax �!��p��A"�XQC��A�A>}�j��u],�MV��\yK�Z^�ԧ����y��E��K'�a#m��b��8����utn2�s�~��>΂�pKe�1��Hܢ�1xA����]0�ӈ�ҵ���D���?��E�v/����d�^��(�:��,6������|�1��ÏL6h�h,��~��ג|���F�ܱ T~�.��c���}j�z�է@��6��� �~��U{:և8����l�0��]���x�[��6
�s�(>\FPm�x��l����9˶5>��ѻ��k��b�dz��xij�	2
�Tw�j�J1\(q <���{�/�鷠�S�~7�S��1��e2�0�����{���$�������J��i�5X��oI���������/�}X��c7�&�����e�mI�NR��U�vF���*t�T,��M�KUyU�+>����C[��4���!���3�
��s�!����[�*�D3��j���:���I�]�o���B^�7nH���ʞ�Y����ߋN�N�i�y�x�M-���Gz)��J���JlO"��c`��,�����A�`l��y1���^j��؇z2�)�ҥ㟜�k�*y�vV����I73��t��	W�|��\�oD*#��Zָ&�ቿ|Ԫ���$��� �%����lF}��	Ţ��:�E�$:?}ޙJC��b�Ė����=F��~}��Ê_Dh�������uO����s��4ll4<d3
Z�_t�(	���x.�q�A�gGq�l-��U<
���,�`��������8�H?".ޅ�zi��%�~���/j���1�M&_B=�4�^�<H�O�c�w�$���(Ӡ)+��zYph���
X���N� ^���;L����)�ٖ1n��T���.tҜ�?`��g��2���䌥vb�i<�Bs9�*��ݗ�vm�pm�L���ݰ2�N��vI�y�84]���T��|�q2(N��G`��N�;|�Lm%�}��X��w���L�Zdo����R=���&���'>O0Y1��&���|�aҦ�7-[p[y�����O�s�ٿ����!)��B�NM�5�c �k�b��ݗD�cE	S�L�U?K[����Ug����d�ՙ�6�N��4om�V�JC`�o������j�0O�4L�+abj�<��#%Dl�>Z�l��n�"9��DYչq��~�M�E���~��B,j��Ɏҳ2�K9��_va�4��`�ǩ䲦y$9��� 7:<���!ڀ�2��< �����6�?	n�?��<FC�4)5m��a�5��^�E|�됯c��b�������P�� 4o_xߢ���.���P=(\��jBe�|�ꓵ�����������'�^7��S��9V�Ƨ7!wjKK��!t�+HȺH�U�Ȁr�!0p�?�e����Z�t�l("�~6��v���J\L�ҙ1�{}��%P�	 ?
PF�jn�e�^�g� �1|�Ii7E��TSOꝵ�Gn�W��/�
����$7���z!v���)-��&���+:$ҭ��]�UL�o�^��QGr�F%�2A�� 6�Q�nW9�_&֘M�U�bN�;�-*Uǐ�k�TFB��s���#ޭ�w;k�� ��a�H�����M��D[��9_�92&XD(�]�����VVR����̃��[�,1��xw瘣�^������%z&��fX	kP+zQcZZQs{��t�����3�B2��Ń�B�4zr�|Y�}�4���k��il�]�e��%A�o���8=�v��X����e�]С����Z����lpش96�C�bv�X�)�kPp2����O(�k��8H̸25��_�T�̜�ƟkuUo��Ql`/�\9�E>��^N��t�)���"�CG�+iGl>gL�Z� X����#Yϫ-��pq�f��f��ǋ�~��j+E�7D<�%}j"�گ��֝1{!�P7#����8N��\TP1wۅ��A��A�5oA���8'��d Lr�@F1����K��Z/{GM��z�(H��@0���*Ϡ�t��ޛ$N�J��/ϗ�2��Jl���F�8�%^�Pr�d��9I(Q6>�!��7�!G���)��1}���7��	��z9�1	�l=�Z��w�в���r
���Ì\�/�~���R��7�*�1��ש�G�LIE���ɡ*|�	5:��|jU6�Y8Bqk������&`���sr�,�e�]u�O���/\S!;_�a����Ӊ��R��Xv��o3�T��I�yb$b��<��W+�����F\�_I����
��/�a2�(Jv��3�f�I�+�b�6?�:�Oǽ���I�Nb.�S�x����D_�ÿձ��=Qx�Z�=�?�g<v��D��Ȕ��~�*�~�9�7�R�?O47����ev�����	�f���Vá�F�[���^|ڻ�(y�&w'|��̬0�s~ރF��k�����������v�Ѓ�p����M�ɓ��$�����B�zg��an������G��x;�)�.��u���Qq?a�E}`u�0��"VJ%���.���B7�̼�h�����	iu�>���DK���F�U��5�!g��~CNg�gk&?{8J���.3�l+DL��b�K?ی`?"b�D� 8oA[�K>m"i������T�-
@��[��$ ��+�26B��vB]
g��26���VuYaPj�eS�5:�GR�����X�|4J�-�Lw@T����+�ʱ�t�_B8��Ɇ�l���)<����D8<�cΫ�F�GZF^K>��;����V�g���Y�%����v����V\�c��dD2�,����/��B�5��e�żGf��%�![+0o`�?q�����#7�ZTP~1�g�PTv�uC'<\XGGOmQ�w�r��7Ѹ�
u�5�28��B:��I�r��:�ߑ� ���t���K�|������Ѳg�n�p� �F[�������9\��Tn�>҆�\5HY�K@�N�oBV���>)#W��m�x��K�IPE�e4�̧a8��'��
�;4bK/^�0�R�>����_ȅ;7Mn�Zw ʖ���G��m� ���9����{�f��'�L$���"���jB9z"`�ے�?�k������Û��in�/u��6�AFߘ�2�_�h�s���w#��"mc��m�/���6�o�tAp.[nS���p�n��x�2�&G-n+�F9�c�<�j5�I�0�P�~s��	�sC���%:�b��W�7k^D<�*~22��m,E�2=�L�b��[�H���B�<�I��c%�x���n�T3__7����X��Ӣee����X�U�V��OpÚ���ar�lc�謼\���c���n�!��J4�@��Z��2t���� &T[���	�e��cZ����i�n�� �"�s>!��'���>|��8k�6Hi��݇m�9囵jn��QU�����~�9���
� �>�'�>��]x��,m�fr��?72��m٥�v7�3��`4̉�;Q�>���5�/T=iƭ��m*�JǦ  ��	��~��"�����H@��V_m}�����w�U2|����f~is�;/<���B�R}��b8�s� I'��=���0'�c�O[��R��W�����R�V��ܡ[�<QQ�'�wG�VY�E�)��M�7z�`U[E�ܯX��А����2���fQ��t]��m�� o1������f�,���6),&��E�Ju��m�������j�w���ȩ���)K�^$Q��@�� �d��@0#��({O���W�n݆K��L�������0����^A6�1�Vj��䴭l��'�#��d��a�9 ]���$&��Ѩ�{ʗ �J[��2v���o�f�7
ӛ�\?�m��E���~9�7i�q����n�E�&G�/A*��nي��sv7�#��������׉'@_��mQ��h�s�>�f�\Aq�L��k0�OuZ
�m3��3 L��۵��$�ò�⧭���|&��ω���Ğнn�ĝ���v!8���v�D=T#p����7��1֜��G8TF0	��Ы[]C��z8ޡ���V33�srx]%A��d�߿Zج���\���t�7'4G�_Z0�w�e8�!��$u�Z_5�H-]G��=�>ZIT�ԕi���봞3^q���n������8ӻ�HΤ䛤�b�422L5��*[GO�_8(S�i�`�l��+%'���N�� ̟X?U�d�D��.��؈�}�A,!�Z��ΒAP~R���-;�92D�'���I����>���4g��EG�If�ֺZ@h�����Z�-y�Ro�$�y<�r�b�9s
J[A����IRoXI�x|��q6�� ���,�@��h��2�O$/����������@8k6j�O[-�*vt��H �,��h�٪`v>z��A�R����#��U���"�(���ϋ�s��+�zd����f(F�g'����Ҫ�
�3s>�5�_A�"4��"���QS�S \q�#D��e_�롁>��Pa�@�s��A�<���V���xJa�7��񰇞�mq�GE�x/�5H�R��D��RǊQCKg���h(���8�W+��w!(���%	�}�p��U��&�o�&LO5׾#fk] �V�����T1���!W���e��l�ԅ���X˟�6o�Z|��O��g���f���4��Ff���ӗ�I6� �����iu�XB�;��	��[���5�*�xn) �дv�9O
��D���*y��7������F����1��i���H4=���>X�DD�K�N	���%�"�ڿ�Qg�*�10�&���<���=�72^2<�%��_@X�q�������8Y�l�u�#1/���&:g�t���}�%ڌ6��]p).�(I/|�C���IQ��"����J�\�voR
�h�v���T1GZ<�������M]��2lj�C$(��|=Bڲ�0_ ��;�,nr�Ь�5����9ܷ��ٱ�(@�?%I�s�:k#�*���������r������\cNU�ofbe	j;�r`܃_�X0�[�T���1տ�Oi���G���ܦ�a��_��j�+�=�T�Q��8o�-s�2gBj��;G�hxG��S,��K���-��V6�g"Q3�6���f%��=Ro�t�RL��-@w_#F��4yμԙ�R���m����r�P_h�p��@����[�ڃ/�&򴂹҂��
�@�#�=���.F{�8+@�>$���<��2�\>-[7�i��5�� ����w�2�w�g��!�}�ʞ�a��6}3�w�>�_6Β�|2�x~����aN��r���Q�5���Kaw�idn;N<GY��$?l����������)�ޑnKY`�6�&È�ځ#+E����0�5��b;ٚ6V����>��Ɣ��)��y�I��bbS���!;�������L��U�T����205'oMl��!^��j~&7���ka�Z��r����B�WZ�H���A)�㛺���3_ٶ޹��.+�2|-ŝ�9�f���q;�!Aq`	��	�<�Jf��l?��{���FW�!�3N�@
�]~�!ې�m���`�س���������k]	�ȏ/�H̶�t��Lmn�$'����
�&�ω3�Iwr	�ӏ�Y��V9��3�^��/\�8ar��c�;�=�7�!73ͽ�j>CM��wJ0�A��1��Ka;)�E��*�cY�VĶ���t�s�l,��e�ڜ-
n�R��z2�����&�C��O���I�
b�*8��z�����jI	9�2�������^:;���� 4�-]t�-���~ݗ���="c����/N�$#v�p��)��d1�ʪ�̭8-�y�W]�z��M?�<���2d>1��q�Z�YYNy��S�2*�+�m{S�&Q�hI��W�rX��ľ:gO��ź8Lس4��jqj"L��W��$`����}��	߲R�FPl��E����<��%Ҟ��s�J�k`';��R�����^U"h1�2rP>Y�]������DYSa�08��������um(JC�Z��Cq�Q�x��L�d�#�`
S�k�&�"Q�d�3g���Ԣ��@�&[X���qG�75�b���+�r��������jm�����p���Q`�2N����0D��������DY�V�6�r�;t�<&vh��X�� ��q�6w`�N�����J��B�iBQFě���~�D��o���w|p�������_Ċ:��TD�$��%#�V���<��h*z%`����)~�m'Mnz���X@�M�eX�8	R!���UO{.�NhE~?����홇�T�kg�ƈ;xZ@����X�j"�]�a���0�_��%<, 0㨘V���V�A��o����(�	a����!�vA��,m�e�Ù�6�}B��S�A��_�(��J�{	}�
��n�]�tX�"������DFR�����L�Z'sgiQ�����)�Cd}�ՎV���S������ū^;��S`����a��o�=�|���ՐZ��vM��9b~ؕ��|����C��| i#����X�a _��w>t�1�Im�� �N��z�^�Р�`��#}l�A6ؽ��5�z��R֏�;ڢ�B��Ʈx������Z��l��k�/�l0�&�0:ʣ�ͩ����Y��{ۇd�o$e���	��0M(*�o#�Dh���"�R\t,�jN�iK��Y�
��ˠ|ї���tD�tv��-B�E�����۩)@@���=�����l;����G
#��������h�oI�ax[_���/���*�v^�]�"՘�`1�������%(�}�Bň�@��ªe4l%$����n;^�tfB]~^�����)s@w�at��L�]��'$���kf�ћؤ䙜aC�j�2��O�:%��|]5�����x!��>�M��S�S@�mfA���.a��@�g�!J0�l�{��TLf����B��s*������bʒݎc�(VV!���7�3e������x��Ʊ�W#�q�Y�۔8����0)b�� ����s�ԹT�%z�f&�<�6v�����A�x7�^�	ȱ:R5i�rϒ�W�'�����+�G_�oBO+��X�RtMM��w\��|�ή�FEc|��x�Q. ��Ʌ;=
��^#I򴢞x�Пe�s#'��۟#_y'����!���{y�+�p�^��w�F�`�pP��<\`c��|��S��~~��Q�<���������:�����>�P���D�w\4���0��*��]�s!6�R5j�d��UI)S̞�����~q֢���ӹ+3�����v�	֫Ǆ�y #�$��|S�*��b2���_�����\�'��s��G�ݯ`���_�Z����=�� �jT8���V\*V��)���z�h�ߥU��&�|0��T�����P����]�|e�1���6��Cá ��$�Bw���	�9h�A$\�ʍx)������WZ�~�NN���] ��� k�d�3��^�a�\��.����h��U�!��rc�h�z���9�&�d>Ŋ��W_����}��LծPO����3��/���c��C�*tL˜�!p?G঑�m������t�;��]������2+o����f��5Ht�I@P�%l|�ǶFJB��Zv�'�Du>̔� �.rX�'�gobH�8�A�)+�	!�+Ͼ~��4�F"a�В"�&<�Բ����KX~%����>I�3�ŔQ���]�z;��e�V
w�]�`�s�0�se �� ��U���<���5���ۑ���z�$���1�@Z���i'E�R�@����s��Aj�y�E���ύԳ]E�.\��mT�g��LG^�Z�H�I ���Ul����)qf���Yǘ&W<�Ϯ���4f\!�u�M����_�;Ky����6�~Px����a��]��զ����D]��'9C]օ��K��ı����#�� *4a!��ӕ� ��1ǐFE�U��G'?���z٤�$?��k�Φ�����X�VؚY�������7�kI~)g��6�_&O��SDތ�+�oV�N��0�%!��=iEpY�-����
>��J$Q�z��l:��-����.��_2�v�I";^髆�^�<>�wY�nX�J��7Q���~]@��ת����&���#J�15�g&2N���ϋ'��H��֞N�B�-3���l�A���ae�7�$�Ed���jr���?/��k'�B����[r��@�´kR�T�l����ge�0�R75鶬�<N�������T��E�R}o����Mq�O�����v�2"Ŝ�_dJ_|����]GD9�}2�P���Y�����ץ�v���(���?���hnҡ�q[;�Hs'R�����@��항�;���@��u�Yi��.'��������] �j>��ʁJ�hN�Ȟ���@DI@T�A��%�)��:�F5bF `��m���G!X{��B�_��5�a?kv�Uq��'٘������W��^v"<8�����X�S��m(m�<t���^�ܱ����Bx�&F��U�$��U�e�s����Gm�q�΢���\��7�2�m$F����7Ma{r��p
*)����h�.�4����#�̋6&�W(�@�YH�{υ~์�J8�������@7�G�"[���˜��z@x���)�*����b����"�0Dɪ�	;u��K��e��uv���0�f	pt��9��ZU��[�5�S��9�7�H$���#��Lb8��x�)��!� X�dܔ�/����	���?�B������o�	��Z��(\��"���y���RM�
�O��GEw���4��)3��:�KŖ��2�.�X5�k: ߕ����I4R��X�2�,��N�}����b�q�`��}����7�*yW��[�C�L�  B(o�>S~���*H1�,бw4���8�7H���y���"qX��b��"���c��s�D����vuw������ͯ^�l�w��dl�+�TH������[�F"0������G�3?G�Z�'g"�	��� M������P�^�W���ENA�9���y��1��C�Q��y� �µ�8�����k$�P�E
T�u�Kak���4����+G:k�$I�ď5�)���i�9�׎������Iag �� �Ig{Ǎ�lth�8 	��X�m�.�ug���W��ּ[w̢sD'�J�}�.�[��P���A��9��9M��ڝ#�#�
�6g���nT%�NGC�_^���dMo���.�Q���VO��V	�pUڢ�)b�?�F��%��n.�*�����_Z��K��t �h�)%z�]�َ�/�=��N�Q�5㦾*�Cpf}C�V�S>F�V��n\v�HR2��φ	+��D[�^�ݢ�n��Z� �;��TN�;&��F�ݝ���	sj۹b�����B��l��Xtc,c��<����_��l���B�"�S@�8�
˾U��dNgJ=��A'A"j	���'� VЮ��Ig�{�ի$���m�3V"�U�����>p�H������ueHeg�^��I��C;d�	�y���,�l1v�k�k
#,B'�7r}(a�]7�Ff�����H]��?���Y���C�׉�9��c�/��˸�����1QA'���a*�=>�W4�9_J��J���5�	�4>�u)�t�9�ٳЉ�EBdH9Y��T?�m���Y�!i�u!�h��ї*�/X���[��)�zk��������i͌�;����9���?�pP4)�Iɏ8ͷ���_d>k19I�m��"y�'��u�ai��E�	����4�o�vI�M�߫go����w�&L��������]j�Qs��ڵ#�]�w��"�C�ס㌌D�\M?r
l��*�ؾ�J�4��ƞ ������:o�sJ�93&�T�T�| �O�5^�f�5���>����qf�[4�>�M�_�c���R9����K^v
�y���0�A���KE���B�d!�=�4��Rk]\o�(�Vl��nx ��Żxe�R^��Q'�o�۱�F�yt��� ��b�H�]wE�M�#kUՀ<��ioH:spč����t xPz���;O�Yzl��wh�ʲ���kn}��x6�&�*Y�Y]�ʸTR��{��Y|-�&lڅ2 V��
"����s�&>�E+9�A���;�K5���Z|����R��>��K�Z�C3���2�Hߠst���G��$#_p�m��W���2����ʳ �&(��%V��]���Ͷ$�]�gD�'^���C�ޕZ̖��H��	�o?�e�NI��#�].T��FK��&��`}��ժc{ً���w�ر�z��SqF�}�}�%��Z��=qQt�P���_������!��f�����|v�
y]����$����-P�y��Ӂ[������4�c�+��!u����n(k��i?�����V/��܉�G��[]X
լI)��rd{��K��KUQ� r�{>W!p�N����x:�,h�}��E4��-�X���E��GF[l|*f��C�"}�` ����w~��Ra���U�;[���R�)(��#����.�p�����;���!O������H~x��9�[�h��F��/�&yМ�$I�h~���9��8�=��jY.㍖x}��.=7ٱv�"w]�x���*���"ܕ�0Wj:iMb��~�0�%yi����4>}�rO����C�����w��+��%�ʾ1������^q����W�֋sIN�f��F#�A�ô�}_��3��{�*��	��B�Z�`�ҵ`� ��E�3������^��=|�}����5i`E�3�l�{9y�o��q^�>,2��o��Z���8� �պs�����F��9���j�wj�iN� C�;3z�J���z�Ck�ǖ�����x��ev�@���u�uq���`�K>
�=4�J���r�"�2`�~�	�S����T�8�>{4�|�rI�H�R�	����Hs	�C���ˣ���?��N���._�� �u/a�4,��^�L�O�y�`1�"�GU{d�hX���Wd��|�Bs�H�ڦ���Ko����ia����HS�䶪d���
iw^C���Ҩ�B���Ew�"W^��I$.E	cǪ���ì��t:p�l��������䯺{��� ���h �a2G��[�sǒl�~AfY
,��準�+־ϲvڮB�~[�d�ǋy\�*���M�����}���C��~h�D� "0>�
�8 Ie`�8������{��w�xp���7^�+�Ĥ:!��F)��.���_�1�T�Z����F�v?���ߝ�������V=M���)�t���>͙�z�/���� 3��8G�W��wv�ç�f�Va8ԛ��|Ӝ �S��t7D�Dp���[��
�������Q�����|Ug.E�D�� 0��3�񨠃����4�0��2�Q�vx7_�O�b��m߿�K�a3�F8�7�`�� Ǡ��Pl�A2��5�MO=#����D��&�$$%���ͱ9CqI+Ø���В��-q|�>�����XD�X:�;Z�$$u�A���}�KKZ�;\��=b����.����,��Pǯ�c�k��XyXDo䯉��v7Uª�at;��v�a`��?�,W�><����We��;g��R�Zt�j}<������p&]Տ7�G�Ɂca]�^9�m�WV�����jԀ:�M���b@˺��e��|��3�6��a�3�ϋ3�\���g�h����v�h�x�5�`�b ���!y�!�҇l�"�S8��L#�`<Q��V���m]����T~Ƹ�"�B=����S����<}��ݪyg�<���]�8�<�u���nc��^��[�d~���Ԭ[�NXm]M� �ν����R;�ُ2 
-5a�I�$P��"x�p٦:�$�ú1rH���LqD��`�D����V���F�q(�inFL�	����A��w�,�A��b��ګ��+6o�������$�NX����v���;y�iؚ(xOH<�J?��<�7����9-�l�?ICVi�S�(�����j�.�#�}1��]F<JʫSE� =�g�y��_r�����ɛR_Qcx*E,�5�AI��"���Y�W�����݊tp���u�{�fS�e���bE.OKa��B�B�g��u��{R�x�Mv�ta�ˁ���>��b}ʟ���C>K�-=���1��Ԥ�|�_2ѾIV.R�8%�9������-�`!բ	(J��b���l�'������K�G~��7*�O]��/G�63�szs_ 5E��g���$���+m�4gr,/��A��9v\7��
�� Qt�J@'ȄN���IwH�1!*_S�A]�5���4�kb��1)��x� ��Ās9Ud����Y���r��ub$����Gָ���*�'m�^�$�t���)���UrN9���e�M�ߠ*"L3�=?����g3 �#)J�E�N�7�&�F@����jTGC�h�*�s�$�7��i�o4W����9 �`>S&��8/;��B }"��:Qoz��_�̌�;�)�*:������z���C"����p��$��ߢ<�"��V/�m�C@cKg6��ḷ�n�7&E�`q5�Ky�y&���V<Щ2ZV[�O�׾�_��Vy�7��?(�� �����*O��l�!�^�IT�}t��V��|0dS�av��SJ��ʅh�b(�2H�S��L�x��5(�mc���|��?�8�Vz2Jp���U5�s�wa�< �vm�`	m�|JkqR|���\�R�I8�ѕ��� �ΠN�����6��,�� *`�n�y�sS��������I�N��T1m�E�e���<�\��:ɏN��c#͡/g�Z���n���]U�-ꋽ�q}�2���%�n�>�S�C����w�{E�q��_E�Yf�h�ᯢ=l�w)��� ��Ѣ<T�I^��&�T����_A��Y�����g��m��x/)���Mi���v�͢QU���HԬ%?n���\J-ЇJ���}tm��3�����ʗ>	���=���T�\'�r�y��
�>nN���`�6������-_`�Ǽ̮����Q�j%��v�����s��,q$�=�3�lҿ�0�n�i���>f�k���9ր|��e϶d��K�q���
o�v���9�ƻ!v�
��t��v{Q���3Y�ի!�e���j���¤i�x�/џGwo�w�����Q�c���6_||��P=²�L�	 A`��y�07�� �,Iy�֔g`{Cd8�vJ=l�k�]��B�.�긞�3�6!rLU��jk�����h|�lu]�C����"�O�_�Z�+иb�p��VK�� ����T �����w�i4���щ]7���J�5c���GWnn_�]�N���-�c����ƿ�D�_� ��'�9y5�7z�7��1�o(S<�s����7���/pwMw�<
u�(��`z;I!�E�ӽ�^��b�a�m��'c+�EL:�Aǿ0�k��!�_m]�� ���C�r7mцʭA6i���j�eB$| ������inyqs�RW���o��a�|閝����Axp�G!�9A�ʮ)���a�&*��Xw])cR�����P�cPEV�'�Ju�{��pB.{��g�JK&yM0k~r�V�Ss�8��o6�ծ|���b�q�A�Ü�i4]�;:jT	����9�.>�@�qkэ+#	7���]4����X����+��1�U�'�ۏ��>�0�*�c��v����u�Ǩ�2�fO����z[۾;��b�~�Y��r��˂b����������.4u�p��(�Y�,�u��Qޭ!>�֫nF��tA�o_աRc�ӗ���c7�ev�'�/�ः���A��|!Ȼ��S�V��6�O��o�C�a��n(;�������+V�`\vͽ��n�޷72=ĲX���d!�!jd)�JN�!���N�����F1��M��wm-Y��m�V��3댆�e���?��'�w�,pٔ��;DP}�΍��U��
���o mҥ�Nu`(������������D\˻0tt�N��Xŗ�Lx2�!��I�w��E}��S���q�{��=�~;��� )�����A�LW`ū&��q�M}QaV0��Vʰ;~#�����8JO6V����q�>U�=�"����h���i)On&Ĕ��9+h>Q'�/V�n�I��{�&����[��3#n��_�Ǽ��8 s�)��@���S����>��M�� �7�s�y���_�nY �櫥3g�É������ż��i�\Mz7��`uK!�ۨ����N� H����F0[E�g8�I�6�!/��$��N0��E�n�@�*(YaW���`B첵�&l�ak3�x)0]];&�e����a���9&M��u	$���Z��`'������z(��%�J�/��z8
��	j�����Ԝɝ�~P&���@Ә:�nb}i�*� W�u�?k%ei����?�R�(�CI��u�G*����z �����A�\f�f
�DN��P�\׽ᩇ����iE�f����LK���؊I��/�Q��=Gg�Jۀ��x j󯡈5	^S�דT��Z џ`ᮓ�'���4�6����I��aj�5%k��8�S"JD��m"#�����5d�]P��#��<etw�����̓U��M1�X�Q�y�� �����$���T�J�e@�*T�(�Rav&+�
D��FܙB�ή�����VT
��A�ׅ������|wc���9t�Qjb����rS��G���-�4�?��zaH}�D���d?��@�ζ�_`�~��@�}�4��5��z}��P�H�X)`p�c����%��%�n�!6c�K����F�m�_/��r+�:I-~J�W��	�6�;�ү���C�qɝ�~'z	λ �&������#��3��������kb����������o[�"�h Cw5�sQ�R��_נ�=7</$!���<KL��jȓ�#�E��$P2��H�#gM Mz�0��ܜ�+��^D{zA���9��5�i�z�=!����v'�[KҎ�Z�0��$�G���<�DϺ�.�+�j}�?S��t�i�b�>�p4��Tk�6������A%J�G\�rU}�2&�h1��8��w������Ϻ4|Ya��R{lR�(����I�d���so '�_�׋(�%\�J�o��d\ꕁd��׸�x�p�Oz�O��ެ���we�ۡ_\�`��#��z�@� �T��?�mL_�
0&�~s,�kӄV�,�R)IG*O����w����Q�m�
��r��$r�&�������e<�ڸ�5���Uo��b��B�w��4#�v��˶�Yg6�d�<�]��"��\R���z|�=�f���p�\�\d����7ϴR?���gʌ�P0�Ի�k�����
��'y#(p��,؄��`��i�(Y�/K��4�md��yb�?q�a��躜֣�\vt������_ ����G0 ���C�"<+8'�Tc�R���fVg���Z�@6�[�iܦ��wݬ�7���;���7��ꯜ���W������k#�\
U�?d�R'S~����
:�׼���:��"����D~I
�ɞ}���!>����Gi�i�L���g+�[M!�!ۄw�N�KA�~��\��m�������[��_}�~?ǖ�x.*����ub���YD���2�d�R��@��C����)OS[��L} �!�W�Gt�ӣg�n�:ì�Y���8<����̀Q�������wa�A�$V1'׎9ͩڙG�4���` t��*��)X�uR�3������+��疁�z��O�#K� L[�e��Q}����d}�+�K�+�s�W��b��h�'Py�6�C�{h�)�2�J���=�����������s�!̎�#9��ϊC�ӟ?I��sK���ɭ�{D��q��{LYC���d��aH5�O��n�T/b�25�6/R�<$�egV��Wܜ|<�*_��ꄉH+�P����PH y�[�	�����ªU�g�	��U� 7x��T2K�X�j-��UV�p��k�;�\d�}!�yR�'nM��+^�K}W�K���QXnX�V,�I�^�R�^��I��M����IK��4�	����c���{�3DaT��a���^!͍��83�X���E��>o#j�p�bR��`5�UCൣ�U޼�����p�@׼���ݫ^�LT3:�3W[�0Lѭ�%-͉�����~\�41n�oGJ�x�����w5��"�Z�ģT�����{>�����S>Ck�-�o�b���KD��d���^�/v*5����&X�v���.�w\�Ћ����2��#�(z�#��: $ҭ��.�,5�� 눭��p#f|�d�0"A��)���V��t�Y@~�b !$��`��r3"p���� P��������D��¥��Z˦+�<��@�C/��AtdE��a�%�t�� �<���p/=Ƕ�K2r��b�A���g�h����+�I�O5������Jm�k-p����%���e����Ǚ%�Ūf~y�%��~���K�jVʤ��� �OH����d��gFc�^:U]J$�ϯ�p�՗~��a����MZZ���~�P�����d�àIG���u���xO �/q�O�:ER;��ej�(���bLX�q�Ut����~G3�vh��4v��o�����5�P��ͽ�5��X{����@a�(�w��S�k��2[t���~����/�#�G��� O떬X{�������	����%�/�.pU�|��)���`�X܅�Ga�^.$RnYl���8h{	�r�������/q���3���**� ����t��B�;+V��M�g��{v���AFv��ڳ��G�����IB~	�_��/�D�&�,�ގ�Q����w0��r�S�0��R�7��b����-�����%�<K"e�m�L���a���E�w(f�D���ff}X�� ���*�8����w��rQ��z�L�����n��]ADf(8�d��LwZ��1�P�7]��*�cw�\�2�ǐ�3�	�«%��0��O$�7,�K�S���@\��`�3f�$�Fim�U��ݵk{;�u'PT�-��F��i�p��=�����'?�ǵ�O}Լ>6�b뵋!�09u�O���v�}�!��
|kK���s3*�8X`peb{�]�?6����S���8/���8�5[+����z��u�h��j7þ����#k��C�]��MLr�_�"A�(��K���2�l��Jk�3�+�uE}W��1龍 I3�=Y�F��b��i_O �0`��Pv�LBV������ �}�M��|��Q-}�FN 0�v��;��r��[�k�3�Բ"i��{�
�4�M��'���萜f�����g]A֮7�'�b��,��0��[�bv�խ��6G1�$\o�Q��w�ȕ�FT���8����	/��i��05<�U�)%;�T�gKB
��>��J o:Y�Q���c�R��� 秤o��ǳ��0�qzgvB�d�P|���c4d��L�7�S�,b��;#�҈$��c,3c�����
��J9�S�ɲ�U��fvw��B��G"��uV��2���GwQ�x�O/����\��6I0�Թ��G�N?{�!��7ۘ~�33zU�'�<���/|F�<��/�_�]/�P�oų/L��?�]7M����ц�Y�w"V���q�q�nt(��EK� �G�O,�^�D+|��bH˺<�,���+F�]�^Ȍ~���6!�m�?�ϯؿ�APc&P?����e{Tp��Ǩ7��U�PST�]�T��&����ݹ�t��I��C�q������9�@���}$���v`q ��;M��̷8�.,��	��@��'�~d��9#��xB�ZC�#�75]���}�Io�{8��R�8 $yz�+~���� �s����T{����� D��!YL�ފ�ú�;!��Zzl�ʷ��LO}W�/�s���V����#�4�)�:���C�-*M?!�Yʗ�*�+j�U�eT��p	�T�3m��c�� T���_�o\t��%Yٻ��%��tl��K��n1 
0�R�,�Y�
K�0���0���~u.�@#c� �"�A/3a���Ka�������gG�V�p�(�f'z���Q[�%%�-}����*e�Iĺ ŷ�C�=J�uL����&i�����⏽����M�*��ZF���o��b2k�k��S���D�)�w'ڛ3��a�$,���rf�rʍP/p��Xk{�ά����}`8�7�z���.�S|��`Pf���ZI�����A�Ab님
�h��w�����7 5'+V.�tp�A�g�3��^LFǧ�Y�MB�:�'��3N���OS_i2Olv�І����ه6�C������%.��(֎�0���qՑT��l�}B�h�
���� 1�{s��-(�\��T�exY�S"���v�['ihe��@
�R)C�Qik���罚
jC�������a��jw��FT��X5��O�i�� �=�,�#�O��R�9<��~rVQ���M7���5�Շ�V�&��L:�|&�?�	$בy*�{�@%�o�����X�T��ҏe�u����B��K&��"`�}"��N��h���oԶ�/�-
7�ԸX����˿]�@���q8^�}��T�-n��~x�,3��(�q�K��c`4������la4Ή��m��=��ٹ��0R�B�-���{����¹�	\��Rw"#��A�K���ש*�wĹHc�!�#ߝ��Z;H�Ď�Y6��ĩ-����ȹg�^����@8�s��V���bL�BF�t�<k����$�'Jv�p@��k�G��oE!���:
v�-�ַ9r.�����6�:G��z�h�l��R�	ͨ�=+Ԯ%�� \�5�UD4̖"B���B/����XP�����5��T��'�$�f�J5'im�$�%�$��3\���9��ޒ3N���l�0�f\�r$&��)֯5�Vz60ܥ���&^j�T����H	f&0'��4�Cyե.
I�PqTr"��L������7���܁�w]h�;B��غ���2�t�
@ʇH�v�\�x�@�G���Z����9���q���*�{v��Z�Lo��C�IH-Y�8��@=���a���K����Uu��s�.�J��Z&)?Miy)�y��Į����fY����I�� �`��&�MV{<Y�K_mI���*���1�X�Z�\v�h1�v�v��O�Y��z�����n��0�e`�����CG ��D�t+�Rg�w��a��S��d�Dh��AT��t�1Q>���k̝&^�|��T�~J<�.�v�x���<G��;�¿��+շ5z)p�B�I�Q����ʮ�-x�r�_ �1h�}#Y�K&\>�p�d\�<��Ti��g���f�J�0������*�Q�VX(��\�iQ_>�ႤE�/��i����0�]��\���⾸��p���L���
7m��8�ۙ���H#��)�m���m ��S�bL�V>�$���! ��"pPb�뮖�>�-eܮU߿���x����08P�]z=*�yR�ƠPѵzJ�����eס1����ބ~���+S.�*J+��a=�w�]j�aR�?|�������h �Kֳt촃�9�����No�R~GA��㒛0�"cN៫�S�VI'�ݣdT�z�
H'JA'�9.	ri��R>�`[���'[�w�/A1��U�)�es��j��	v�	\`h�^���U!8,9���c�e�o�c��b���(N�~��1ldAL\������gP�y�ja@�F�}}>�VN5�T5�CŃ�d)Ul3��
�/�ʑ�
�>H��T����etC8�ofE��W5V��z0Y=�RR �g!w󀂁77���ŗ-�HK
�j�n�B�L쑣X��!`�������m�}*��:O&�*qU�4}�F/p�$���G�N�o*U���,v�Qri�5������.1n�`��Ѭ�>�h�89߰X�R;N�ܽ۵Fȡ��)۳{x���TA�!@J��ӷ�n��7d�^���@�����&�P��d'0
\ �0�� 6�Nù;w�kjd��J	�"Ym�f�.����-)N�{ @l>d0U��5�Y4(�������6-��s��0>OO�X����cE�
{[�z8�;�>N5���=�����]'��p?zx֦F�p�]����vTK���/��LIy�i)���l��uT&�[�>3Vˌ�IK41�a�׎wŌ��q��a�����%�ÀՑ-�ZM0�����t����Zg�Q!�A5�� ��+>�%+���(�nu��c�Yo���	�~��,��
�����n^�x�beЎT����.<�e��0d�!�=޽H&6� cZW\����*��E�%E9柜'	�i�ץR��ږ@ȿ��q���)�K�l&���6O��c/(�g �+�~%��:����X��%��s1�h���T;_�A��I<�V����2LJ3��{Qc��i#H��̣9/�#�GDg��CJ����0\�#��e7��+�/���C�>�j�9�$����Ae;��H��_�v��L$x��S�x�f���*#�BR�b�iiJ��H�jht��/6�y��$�bvLo�EM^#�7HLƭ&֓dy<2܊MH�_j�4���}�|B�@�G��Z�We���0 s���6�ANxq����!���V5�����gS�D�2Z �XcB��5��Nn�0B��jZT�t�~�/����(E�Ks��v�oI4Ui���gM��N"x�ds�5���K-����	.���6'�^ZO1]Rq�j*���I2�. 7���Q��7$�/~q�0��!K�Soz�+T�̝窆s��Y?dꔆ�F�rCz/3ato�>����$�V�U	ѣ�k������}���<�i��K�8���L<�8Q�F���7�6M���?2�o������ו�p�r\I �A����[7��V^�VX���kr�:eNk�!��f��� y���^Q��u�7ܓ�k2A�w��&,���(���Ӥ�R:�vЌ��h,R�tȹW'D<]2�Y)��˽���K�X�M��`�\��Ѡ:�k�_�D��ۄ$����ф�$�|\�0{3��	bY~k���͖S���I�8�%��[�d~,WR��[m �應f3˹=d�%��&�0���n�䦜��i{����w�V>m#�_�ѵ�B��ݚ	��������cLf�B9oh7�V�
��=���ƕ�4��T�C�%l�C������A�M(�4�3��*|��ZDg������0��n/���i��MH�ӭl�ـ6%����z�XyD��~ibr���:.ݷ7���<3z30��Vd)��R��5%|-�UDA*Ӥ�\���iM��?&bP����QwW�ˑ� [<���A߰���}�[oҹ�=08y����!�Z;U�Gp��y�X��U�|󡉺;��I�1e�'!����)8u�q##���d(.6��Ь�bn���6�g���4��V3N���9d�;L2���v{�?�o"����^�X=t-���\��?��_�� � ���^^��C�b(��#VB�1h�"9h��ެ���&�I���"�&1���։���H��mC4�=���`��N	Ծ-?�r���t�>%��v[یz�dWņ�<Lb-�_��<�yhP�߱(2c�R�7�f�M"i�L��������9ֽ;:C"O&��&k���T��w�����gh�wA2~�"3�d�*�`�7FU� ��63���B���!��9!\�Uăs�>�\��/:#6��D���X���p�NuA������3�\�mu��B$`�؍}!L����#V���&Ǵ&����@��j����,}�˙�6%�06�6��Ǧ%R�gƀ�>>�\�Y-�8FX����t̓��������r��|í�k4�g��[��_�͒m��l�f�&f,k�4��f+�E.�Z�_�%&�j�q�._�I� �qqr��#��n3�h�b�ߖf�%G�Xi��r���Nl�/�h^�t�$�GO��Q��]�b�{�e�?�Bp�jm��c怶�1���jqY ��"RT8�GX��@�x�F�����m?N	TB1jU��5)�ϖ������w��`C";p�1y���Eժ��T�y#�H��%�L��Cvf�Ѭ~��`I���k�ɫ+A�2|��D�2}����,��BG�lC�J�>᳏�wg]�����$�"'(�SG�pC����X��ڲi�S&�e��Kh�&��o8n`�C|Y�oxP��<��}�|�a\��~�!�ߝ�z�T]٩f7_��!to-�1y!��b�1�F*Lw�Z"F��d�eHFֈ��2�HC�ʱ͵�3e]��A���:}�}�כ��j�zgZZ��WS�U\�@�yoKC5w�z��g��o�|6����hM�Z�/�����tDN�s��D~��ά^�����=���#]�mS��*��(�	6�ch�b���6_w�`��τ�O5���46jHْAn0냻6j�k�9�J�G�I#��F���U=�Kr�\�ؾ�&���ܞ�0w��51�NhJZXN+�@}�̜��430�d�h��H�`L�4��G��o4���酨i���N`�?�N��F
06\�	�Y��h�p�7��~	��ċ���kJ#v��Uj�s�@�OW@�UD�y
h�מd#D8�G��&��1�:?qp�ZS`$���kw�f��%#�+7ED�<-�ߋ���m��Y_��<{�x��S�pe�=�O�~�MA.u#l�".
ņ܌�>"��q�U �]j�G_���L�.qs�T���.��IlZw�+����qB�
D���6ș������AB׺ya��5���kreM�����nqcl�7^մ���j	B�������F��SyZ?!����u�����>ޘ���A��<��V���>��l����e?,���K�y�(;���M҆w_=Ȕ�{$��J<�ܩP86��!�hŔ�t��u���k5=C�����BŅ���Џ"��#��O����؋Y�Q��&����τ/L���?�'���o���"^=؍�%��d#��:�t���޿X�D�dl�ӟ��J��GM^��lR(�*!�5�, �1���)V/zGG��d<嚚h4'�ﭞ��+�������'��M�\��
�#�������p1�z��oyyT��N��:1ё���}$��q��7�e~l#���o`;;{ᩆu5;Y��'%K��F�}ή~�����Q�ǯ��l�J���h-�}�X�>ĩ `gq�z�tv�Œ�סv��,�0cg&7L<_Yӽǧ�/2�b�G�8�]�9IS<�c@��`�E�99!T7>���p� ���o���-���YG�x�R&A>:�kW�#���?9����/��R���9VZc���J��	tF����;��+����лzfȔ�G`��~Y���"����NB 
1T����ˏ�q��N/�Ar�����f�J���m�f�	��tG���&�'�<�\kj=����&n�c 4Ħ���Y�y�x�-���Z��!�	@l����8鱯�*���� [[R;r��f�4�!�\tεH+����E��#)�P--�/����.z��cā������W�#������z�{��%%��ϖ ��0���%j<�
S -ĺ!�]|�W?5$�t �!ǥ���!����$>���r�WeJ*�)��kZf����U�+hkTޞ�J��P�d��R3-��A�~�}�!{��x�2|�d�?��
x��l�@q��:I�^z�-�h~i�<���$���M�p��j�]����m�
Q`�a7?�rO�U��(��xaG�*�g+d°�n\��F�9i��v�3�[w��Gf ���z�&E����~u��'�Bh�p2�s��U��+*�k7�#F;p���f�s��q-ϫ肱l�JS�!瑵��+�"V��^���4�;=]�ij��"覧h��%W�x�����ρ��*<�C�ǜP�o�9�T�4O3���A{8W�%P^����y<�� ��i@5 |[�ʸ�� �_df��\	=	F��oF���ό~Ќ��`��ORݞ�����s`V��&P��M��i���Ne�w�����ɪ{���JT�&�g��e�)����<��JV]�a�؎d�z��S+EY�y�ʬ�?Iۅ���R����4_8,��A���H`_�MD�RR?騧98e��.���O�֖����'�6,����F>��]s�ڬ��	Bl���I���\��
%^�u�xe�~�F���4�{ӵZ�췩j��]<K�y��x˘[��DlM�#�G��F3�E�&6��hZ��y*�$���9u<j~}̻�ј��ʖ6�
� �Զ����ڇ�Mo3�7:��d��Է\�JC�v���C�5u�Yo�NӃ��ɗ=�t���m���:�q�06��X�ךR���u��ZR�
_����֛�
�S�Ǝ����}�,����jJ}��U�]�Y@7�"���WC�hg���%]�"�
Hqso�m����F1��@�)7+{��\8'j�8�Jb<��oT.��Tv�*_f,�<G=׿Ԑ����V��]���qɩx�"��r�]LB���I��^��n#�Q�8�|�Bib#�X3�-@������
��H�Hi0�S������'��=�p���<�KҕVrv�z.��D3ɏA����Y-�+E�z�V$�je�����?%Ml��v�/�o�y��1�?�oN���|��D�����������B�P�C2��K9�?$�n�{ l&��u�l)��J�^X��Y�߯�8�;*��Й��o��UAH��9A��q|Sh��Bɼ�7�ۀ�]�נU��*l�$OC^tڬ����Y�.Jqx�nL����0�/u��m�K����c�ޫ��b���W���i�<xo�/S[av��y�kNS�����mX��������.s�5׋\��|;肞	YӼ�=��[��~39�1+m�2�ѿ��Ɛ*a��
��5O��6��ך�(Nmd�V``a{���P��)O��VD��ƕ�h�_���,�O��A0�OѸf��a�aL���W+#��� ���p�&�-�B��FdA4�V~R����k'�lR1�I!�r�>,��@�8���٪H�d��f�Z�����sn^aV�@0S����TOwT�t�$A��@�l�!���O�����Z����N���pkF�HǟT�'�TJ*�N��1X���<�7�h\��31guOV�r���U*7�y���'�P�WC#3�_3y>��J �)�	,����	�Ńs�3i�@��gL*�p�zyf(3�Zu[���,D�s�hS~��i2땁Ѓ�.�.&�;�s�s�z���I3��	[_;EB�n�wef�X���W�� ]���U�&*�H���b��rW���
��:2�	v�;WE�ܶ���檁��M���Hs8uKP��bn�%ƒ�\z.W�v����$-�*���
O#%�Q8�R�tJںqh�8 _Z!�x�g<O(���dDh;��׻�2X�ԣ�ykc��$�i��I�`�W����,��%5�V��� �s�/����J��Ł+�@�w����J:�|�N�o��F l�t�����\̷L��a��y��,�$7o2ޢ�Hp�H8y��D:)��.nA8,�П�3�$�sҴ�Qhq�#,$��\k:���c���n�?�-/��$���w���IՌ]1k�f�x������ь�>���O��p������B�J��QH���$1(sEz$�u��-tG�L]�i���`�N�>�+w�,VH��H-�'f+1��FP�C�W�oj2�w����v��9k�B�fֵ��b�72Z�u��'����&F���"��n_����N+T� ��~����;B���uv�>l���J���i&5��$WP#��; ��b�3�(���R���W�xP��;�d����q��Â�o3���sA�%��̒CD{4�;��Xke������F��Ғ�X��S�_�bm�5�#�?�=sc�w�L���:���M�/�-�yxep6�>��&47�d�s3oą4J㢇H�a�3E��/3�@�JC�����I�����:e�dKicvX��>wo���Aa�d��������'���"<�-�K��p��7�sj�ͬ�Xó�&��H�C֝�i6H�����<&xP@�!���ш�����c��j�fD
v��i�a�A��G��&GgHS(mkv
�Fb�	g��F`)7�YQp���^�z�d����1G_զ`;�������e��g��lx�L��,,� P)�'����l�Q�nGi��" G_.��x�$�	�� �*��$�Λ�բQ">�� �xB���	�F"_��u�]�k+W&`k��ͯ��̉�\����K�amw��Aס��.��x�,'�8��W#Iv`9��1�Uz�S��uAG�2;/�AX߅AR��6�4��G�L�(����7��f"�&֧p�y_ˠD�h������s$�QҹP�'ŧ�l'ږ�e���Ư`�y-�j�Dʄ�݁���P�\T�m�����i3�d���=؃V�а:�ܺw῕$��"�߉ǽ�,
��vk��qJ��lx��JX�.��%��.�0ؗ�ñ}�(�AD���%�o8���of]�Cdy�~�7������u�l\�i�m���{#��W�"��3C&������u���wlO�`�$�隖l�ܡ�$k����P5jl���H���PWâ5�R��Q�!X�扭��8���F�l��4Yh�ω�HX~?݅���!zMd�H�H;��=�D�5��ߵ9�*�h��Y��-kh���f"�n��2��z7�JҜM�7����=��>O��X�[�;5��v�R���Rpi%�ށ4N.�ۢ���9r/���"&C�p�9�1z��o�� 6wDoA%P3�����r�QG/
�ݴ��F�6�]Y3�F29| �}E(������ m��π3�㳑���yMJ�#�h�9Ủ'i��Pt@µ+�⪅V3�aMҖ� UI��h�d�1`0<�+�}�rΧ@��A�!��/�=��������nT3I�&"�C	�4V�q�G���{��<����e������r��~��9���#�0C���[5 ��Ӵ�]�*g@A�?!��@ Uȵ��,;+46��˾t�����E;vd�-��dk��E븀����4;�e#j�;�d�.���?�n�@���[���!*�c2)n�3��+qZ�ī�0�����t��o�y�Fo��lDԹ���릨E}B[بv���	�,i�&	k���m ϯ��'z�����	SO"���u3��+7k���V����ɷ%�7-��.(�"���ֿw��Pv�(�s��ގt[< p_����ע>�]}(@W�#rBx��&hT��+�7L��F�g�םW�Pc��$�Z�v�dVdt&إȮ��C ���ǫ{�4��AL���UpU�cpH� �}MǞn|OT��1O�%�穃d`΢Z2���#�*��N���$�����~��[X�9\`T�.���^�/@f��/�5O���Q�>r�F/+{�Y4M��na��b;���d���s�������uo���<�)�.�"�����Q�U*��\���*��Q׶�Dع?����6���սLqiXR*�a�,pj8)�"����W��K������
?L4[u���4�L]�r�q�F��T��x�W����OKu��ѷ��E�j��\�d�IxCl宋�H�t��O	�/��3�?��{|�C�T"(D[��G!��<��bPd�� ���y��o�$�������z2�"�F�t������O� v&�GKΐ�c�g�,�YRAPw�_~.	�޹��s
T�B�Ә�{C���
��c��TPU�i�*�j�9,Au/R�g���qRb��zq��{���r�;u;���
(X,�����ۥDSi��s�ykL���Y�D���
DM��!�U!(Z��{��I��a�	ofU,C	w4�?Ą	
'��9G��^�lr���m�R�����2��A��Z��Y�
��F<5筴<� yZ�׼w�٢��;�0d�%���G�1���������K���nY��&�J�����	5�n�fަ"�]kx^����_}���!����~��j�����9��^o�-�p�a*�%�UJn�\��\�"�i!�ǉI�L���7�H�S�������6�={����|%?�wz��)x%(�6TD�X��mH��Oصa���A�|Zd��h)lq��ߞg�4�^�~�%uo�n�'�PB�\-A�z��,1	�/=l�s�B<�c���e[t�Zz\Kg�:A�7�>�r��-�>Mn��<F���a���V���O^�kk>���|���̐�d]j��I�iWK�D��Y17�J�ۏ��ݦ����+�>�gb�B��uB��=f&��[y��˘uz�u����n�m��{#c��kf��s�g+^�?�"��2X�%r#�kJ�@I� �a�3�G��U-8�!A��(�C��<ߙTH��A�k=a�̗� �64�[OY��p¬y�.t���4K������Zɒ��z��:z�T����x��|$�^ ��bmx����`��턻Н���4��-V�NH}�]����K���'b>��%8Gwd��p�~����ky��c��b5RW���bx����g	.�����gE��T�� ���-7sԢep�&^p�IAE�.\��v���s(���~�nȒ�+TYp��|;�Zp��(��M�'tH1(���!�z���O!EF/�3�4I$"+Y��1�ny����}I���)玗�Y�I&�L�ɩ�SD:e�C��2�o��*:�d�J%�ƹ��D46����������Ӣ/M9���^�:�k�|'a���$]�Ӥ�7S���T܀�,�[L�K&�*&M�a�u��YmjbC �y��[�D��V���it�3q&��5+�%*����5-?��ےPs�;�dQ��N�Q�/4�rx=@Σ]B\�y@4&����M�[�>w��̬�P�	�O������w��1Ʒ��*�\�-l�yg�����x3�W,�gLG�;��PWG*J���tl�ډ�9g P�X���~ɖ��������5�8�f�����6�篧f}o�x&$����h��,���fI��zs�v�����@nd�%��h�/�]_6�� ��;}���H@���Uʗ�������HЇZ�����㭝|<�ix�+�G��՞B�yNjRy3K$��>�?� �?���� ɦ�����
��f�"BL[����J�)�X�cNE�0j��^t��u�4w��.w���WK�c
�B�莍iC��u �]N�KI{�����Q�RS�N�U�w��c��xفVT�~�����S�"�S:&��h�M�y��X;���8�x�s>�6���/��d�o��V�;3�cF F�-��[�۰K(�)��.�������ri����5���[�`j#C���M� *QCoNSB��XK��
=��,A[f>Qً.d�K��q���2R��JUd�=���Y��rU�Υ�_���Z2��*-�zf5�1�6OO����V!����&�X@��A�ձ+�=f��q�c"bH�Nn�?4�LN1%�C% �}�M�3�Ù�sRǂ��WC����A
헰�����\EY�l��6�%x��������u�خ#���pJ6��L#�ѿth^�R`RO��x &�����jr�(�~�7�*nE�/�Z#��mn$��F��rf;.և�ۚ����ت��U�G��c�Is߹�Î؃�mPOTq�g�Va!i�r
����{��>�՘�h�6Ȧ��
d�Uc��p&vI{�h��tf�'C��0@���7L�,z?�Q�U[��>�����oLسw{f�x5�u�b�88	�n= �Ǜ����ܽdY�s�	Y|��f*�P�/5-T2�Fw~���C֫0d�ЮӚ���T�
)�Դ���To���(<Z������\�H�,�F�їC��36��{���8���5ba��_]�_U���wO�y�����>���'�0{4Pf������]�$��Aλ�L#Zx��|q5����м�K�Χݷ]�^K|��a��a��e8EPp�Ȓn�B �6BĖ��<e�LzSe !�M�K��<��W��cz�:=���J@\�E�:,B����\�wu�� Ct���s�����6�Š9��n�]�w��f��E���F��M2�&d����f�Ug�K�YԸ��P������+�I��2����!��s����n��D�{=��_��q�k���g ݾ���r}�K�p��Rة�Qm���n�{1t!._�w�����$������Z���/	����hp(v� H�̈�x'���^I~Lئ�}���Sk�L�q�Q�o�!ZW~��t)h�����Qq�kٍ��a0#��0���7jT#���:r�K64��z;�F|[I���R�y�B�V(�'*��9D�cs��S�6Q�����kfͥ�<s2��N�
�ʡ��ru����p,i�����H���.�3+���q�BY9���a�D�x6*!�����Q<����؎r�茄�p��}@G�ⷱq����I
��������I���� q/���HB�#�o�W�7��t'K������C�#���� Ӣ'N��%Ҧ�޿���5�F�']���Ћ�o�GSs�_����|�%�?\kU��hU��l���{,�`����x]!E�)!C�����:螱?�>��#�?�x��p�{_f���^De�(�,}C8�I���;��F%*⛡�#�r�?���O|��3�3zb����<���� ��S5��:��vb��o���c�Π�j_����#�me|�-��/_��϶'T�X�4����RUe�N-�f|��)P=L{�^�]M�#�6E3�6/o�G�s�-y� Z�_K���J�IHn�I��8�,��PR%2�8����=�o5,IN+K�X?��k�	�C��\Hw���%ͥM�0�z�C�%��
�p�YO��0:h�҃��/�\�	���u?�[
P6��lVg����8y���{����|�\���"��>����M��5�G�5`�<�o{���nzq�B�M89L��yK���yt���:�AXn�TO^a�.��r�.��9��ht�c5&���!����45}s�"5{�ӈF�H�}6����C�Y��oE^<�g���>v���ۂ��GX�	C�?�h�v(�TC���W։�@�5�p��f�G1.����dO��\�&����R�
B�� x����V��S�-m���d��6�<+8D14�U�Hє5x.�Ù����]�����"
���g:y�{�v��A�5�IJ�`[���&�0&��!I6$�R^43�;/�e��&s�uln���h��ۋf���J��/� \v^�&��o����"N�����<�3ϴ��HW�sD���] �~m��i��SW���S�Wy��%5�%�ƶѷ��ϟ�v���-�I�1DZ=Ḣ��J���*G�$�d�Xt�V�!p��N�A��(�f�g�/bA=j �9�������@�t9!� !h��p������8X�|����Sr	J�_
���#d��p���/��# 9T ���-��~�T��Y�:�J9���G��>UYF�}�!�J�ǉ�SW��F�7���m�kt��"�� ��/2���~&��aZrܺo�����D�qU����@z�ފ�w�[��q�:����=ػ��oߒ��(���t����Y$U��?z��w�s����Hk��S���S�@��_s
�z=w��Ķ=�b��Zf��|�dV���"W���ͯ�#�r\OnF�XB����:H��.�-{d)�_
�@�<m��f���{�/�k���M�Ư~���,)�V�� e�$I��k4Tf��
li�s�|���w�Z!��j�9�pZ��E��a�X�+�9�p�}w�ddٯ��M�J�w(�t�u�Z�"������
,?|�Р���r ��h�4[�K���ɝ���Ac�F1���3�k�/ � W>j��"����7Q�_! g�z�a�u�kD���A���o��{��l	6� Kw���p쩛�]��8� G����'O*�D��Oa��T��`�l�l��]�~��|��;!;G�����0�w�\�?��u>����	m"��Ћ�����8������b�Y��r}��O%ϫ۽�A� (�z���E7��+=Y����F����m��з�}�"I���l�r<V~ʌGF�i��-��ʾ�?�}��W�jc���
�,�nb��L����t���9�H�o���',�ය5k�e�OdVz���3�,�s^G�(�6t�q���vb]���z��3�W{?��ʼ[�0M5�ʝS��2~�ǉ�I����0u�Lu�G�g�7���e��S���vޏ�L���P>.��ao�s,�	9���Rg;8N)����_����NC�o^��rNf��-�!�Nm��U��P�׷����Z�6K�)%g��m
t,�r�NƔ��6aR^K@�#�h)�J֩M�,��i���h���>&�u�y%�.�#'�q��է��/���ͩV���Ŗ��Z�o�Je�G�63?�)D��U.�a)Uc�%n/�<=O^5�^#�/���;` �	�!V���}�f��(P'K�p��R}4048sf��o܌&)V����q0��~��*��I���j97P8J���tM����೦����J�ߜ���ձM �AJT%�y���:;�!"��IJ�f�ى�'"��ԝku�π�:��/���!�>E�WҪKa�}p6|� y����e�����~�ǳ��8�+e����&PdD}�z��M��:T�ȏ���s�C�pk�#��&�(]�	�M�7�>���U��b��%.��em�����`�4�7@Մ�f��vXX��$<�;W�� ��Bz��c�O�D�w�5��ɍ?-�����߈���/~x�2���s�I��+�wM�f='R�6�~1}�Hސc9���ܜS�j�F���'9j�I�	�0�ϻӗ�(˫_�Cv]D��i�odz.���5���\4����]�EK+��%3-��6��-p��N�~��£�z�h#�Fj��$3����R��L���NH���A�MH\Mg�t��va���Ǝ�5�X8K�`�r.Λ-&��t0ޣ�ݣRY�l0�k�O�>7�7��hy�20}�pեR6$2�ޢ���4����I�3��s�a��yN� ����8���<}�h�?: 2!�nͯ8��O��/����j�a.��n8u��-9B�)7+^� ���-��uP�Bh�ߡ�Y�K� ����d�S,����Y7 ȳ����&Ul_��N����sᡀ��qDq���c�:y1"f#G�?�����{�H��t�rm��;�a�B�l2��lt��"��i��XW�S=u�A��&z����V2Dz��__HvxN�8q-�(���XQE�v�ϏL�%������Di*#,hR�K�[>y�1bs�񊰘���N@�aY�(�(쎱<>l`F��Hc����B�������I�hV�����'��	�im-��IA���{��`������i�����[R�D9��FZ[��6_��=fP;���T�C�.�N�)����Rҳ��J�q/��Z��ζk�u� �j?�i�hg[3~�OJLw�,<d��2N�y��E�t���Q�R�������0�	{C���}�1�'ϴB�vc��DX�a�5�R�:i���QwG�"�\U[:������셇[Vl�Z�L��.�C�ԡh�ՎkuMD)X�a�������	���m��&:6C;]=n��P��]�J1풧�q��Xl��ib��@�2�A�E�?R�زc�ԃ�cP)��?@1����$�����ңh勘ǌ�t���o��
䐇m�-K���d�����P�˘~g��`HY���\�8S���瓈�����%j��a���һ�<dL���w��|Fa�� Wp ,���*�!LZ�������kǛ{\����}.
�Ł�J����d`��\���	��Y��#�Z��0�=i�Ӷ}�8�	wg*�U_v*i�Ի}k$v���ȷ*K��W��^(�D�7|7ЪU�6���~r�R�H��yr�Bmv7$qUY�9>+�c����F�d��qE�U'��9Գ�}T[Ϝ���	������|�'���
�"k�-J���C_M<�1���Go��6���U���f���1 �Gk[F�<�Bs��P�VV�D�?h<aj-�j�u��޹�F�E�����Θ�Z!][+�3ьtK��z�d�` О���k�&��R�P�����t�����ZH�-p�b65qׂ������1ZV���gtZ{Ϗq���p����͈g����r�5�R�����e�+,1A*K�R7���}��=k���l6�����M����J��Ň��=',�W	�L!l�d���c��>���I��顸+h��Hds�h"���p/��]b�v�8
! S�@M�KyY�o�����20�-����Ph������D��yg��C�-`�.�!�
��nI�fv��b��J��T�s�-�`�ĵO͓�)��&A�ܜ�HZ���+G���;��h�J-��H
�s@(�v��%���N�q�b	E��8J��Ӛ,v>?���-�Բ"��gWys�hh%�+��̒�~Ϟ�#c~<t���7҃����#J�8������p����c��a� Ml]I^���(k�X�~*���3�������;Hj_ĕ����=Z5����j�١�{���x\�R�"� )Z��"�M���`��-,�SY�͜7��j���|K���䆭 B-�l>hO�SQN�l���@GxrTyJ���p��D��x���6uuկ͍�"H��I����m��c�t��W �ߵ�������T�n�ck�r�L ��e!x��$�r,�l�,�E?!��]��4q17eOV-l�kH��O��WB�I�0���%V`���4t��︠d�,d#���w��V8M
�L��>�qZY��"��e�zl����O�7�(���p��]p%�_ŉH���u:�!Lo�'��`�-g؈S�M .LQI]�||���u�~?���-1��W�^$jN/=	�,�j c��ݹ'?X�g�0'*�bͨ��	��ֶ��a5j2Y���T�K��r�RJ���4�'BU�kK��ϻ/<�2�ǥ��U'�8�d�ٚ��ř�(���sB�9-`�"A�T�lZ,C��]�
��a�䍌")O��K#�����6�q<���2l/�Y�G]tg�xCU5���w$��eI�������uj����Av'qc������Z�i�-D�([�ʎuU�o�u(o|g�"^�C��������=��V��p8���	B[T	�&�(�Y�蝤?��<g"��P)���4p:+��<�N�}��˟8�(��+�.�Vu��A&{�Aς��n&L��lo�5��-�j�*SLT�|�bB3�N���Z��[��])��ii#
��B�ڣSE����%؉:�:��gGw���ɉ�Zz���9�hhO	XZBDЯ��Sg�( �,����/-q�DR!�п��.��	�tkuY3�5������q�|!��
.�3R��xjr}��<�i�p6���!Q�m�frZ"�����(��7Ύ#� QZ�YE�j���Ǹ��I�H�}�~uś�̱y-��S�S��H�M"\��5	�Ue�K�"�"��HV�y���l�}H������k��x�Xm�D,�c���5��EǶ^���z��$����08����Й�*�X@,�*e�P-�Y�>Ze'�Tt�K�O
��5�>��H�<���2�8��Y.V�u�#�����,҄���LzV���1�F'ũ��*��:o��ߟ��<���������DJo�`tL�$x��ҟ��:N}I�:�h�P+ �E�̩|���נ{u�<����l�#���8����c��@vY��K�ۺ�87@̾�a���X$D@����7�1����Cr&��7^��x^�_�k��V$���oo�� [[�D��h�^,T$_�-�����H^,��42�ٖ���:�ŉA���u}Qn@gJ�T9W��������$ e��W.��1�{��	���wD+s��Wq�ƥ�j���H�z�����G{�C����Ħ��18-u�KF�H����O?����̡�V����ŀ�^�/Z]7�,�p�L�:��-�6�� ��PT|��muv�\�{g\� � �w����?Z##�#��0���z���g�0��_�&��`,�w���H��l�VǸ�<�K�枱�@��ӫ�/Q����R7�� ����t�K��=k\�A��̎�6a�x�A-�]L+�u�q��V�-*!��4���Y1Xed��D0��u�w�Fx���{�����׉k^7���s]�
�MvO �[Q�7��<%�@����� v, �
c�����]؆��C�"����Hoie��e\MsCE�F��@v�l�޳Ud��єa�!$��M���S�H`����JW�M&Y�:#]�<��ĻI��K;�k�w��qB�Z�.$`s��L��⡅Ь؜W饬�f^k6��{��1�ݼ���b�|����ڽ�D�f���x���kn�eyq�ǟ0�Z�wt�@d�6ON��]Ɓ�P�M��4J_��I�v�]��LM�f8����Lj�<�S�7�cX' �p��z��M4�������auW��/|h��x=k�#1��,)�$��#�[{�7Xӓ�{ą(�k?#�4s���������#$�������c[3�֌~KL̋D2������ӭy�5�I�`��$h�<�<�������C�P������d)����VL_�x�bt�y��ԧ
9w0Jcl��kJv���;�R�Lɕ�����ʺ�%�QA�=���%zT=Q�&���=��L!5����I�Eޱ�������,�� �ۭ[SM��_�UN�8auJ����n��	�$*�I����+h��V��F6Hc��#�tG�^{P����){@.b�H %j�����yj�g[���N�&"3ˋ��a�I;�n#O��|yr.�F��||+���J`����1�&�z�[�?�w�	�27��r��T���+q2�:��H�X�*�".9�/�$�V��L}�"@��s�����>���S��`��D�
��j>0���o�n;l���������4������߽�)c ��o=�n� RZ��N�V�ѽr�	�? �P�@rHi�}Ohu��� Q�b2^� v>��RPаA�c�,�2Ata��.��s?#1n�S6��y;��X�������{u�[�=8��BF��@)�=e�gXy��Br:�1C�6�P�Ą��.�]�g��%�j,�o6!*H���]�`� �b�xN��{>��v�P��MmFYC�YHv��6�G�\��gQkM�n�Yd61ޛ�	Lj<c~T*,�\�����8k)/�Ѻ���G%����7&kI�Jb�2����D���PήI��1����s<+}�}x9`#�K�Q��!��AU�ʀ|��0�5pS���p�4"��W�Nd�wwQ|ۺsT��&t��|�`^�������r���.L��Qz�:5ps&��0\l1!�qT��r4����ԉr�ۗc�]��m�Ew����)9��Kb�@����8����rEMEB}ʭ�{b�����q]�8�y������'c<S3�Hi�]��n #`�p�8A�.��b}%{wRq��^*�Uq��)�kS{`�	c]���$&E��j��j��̍�D�	բ е�����G��h�	fS���5m?	Z�Z�5OT��������k�_���X�,� ���Oi�hu,v��A��c�݆�ʎ"_��Xr;��7�\� ��(>���%0��/�o#5��J���UP��C4��
+.��Zi�}q��!��¿�L{Q�W8�	��gBu���jA�?��1߹�p�dnI��	w��{����B.)��gU��g�6���&�}�PE�Z��Df+NӰ{��t�xJy=3��z��؀�q��D̛Vf������RN[�*�T�!H��L�1�z �833�@Y����(���J��մd����6�g�lV�o�հ���VD���Hq�nwc���-Gt4�Vt>���[�Hj>`8��%Hay�`v:ۋī��hk�������F�/`4u��XP0
�ꀢ�/V|_8��I�.dJ�r��;��.�3�:D���	�L�}�0�T�6q��<��]V�P�X�"W�wS�����{����BMJ��B1��:z��� 1�W�~�����������lڽT�}6Z�� �.�T]MQݽN��H�RQ����T�9U{�����N�u���s%�|��á�> \�����z���۪ l�Z�3�p� ei�|?�;��&W�&��	�Q���VwN]X�i�T�_���KN���S&�M#ա���vi�S`̓m܉�]�=Ȣ�Rr�~o��)B܁I�5N���1ǆ���=�^P�,ڍ���;,D�P߫�E {6rWRl9�??�������`� ^r�M��ւ��?�uB'p�M4QJ�x�%��H3�#�
Y�*�+p*��C�S�Ts�i�p%K-�ù�,�F��<T,Ӻ����4Imك2�]L��e�+|�G]�� ��ҕ)C"�\?u����S}���j;��G��Q��_Ju�˱����#�	�ZҸ�u��*H�~��A�8�L�|O���aRН�'�IqO[s�,Ѿ}�SZ.�.��pg0p�3�q�ND�"k_X��	���v���`���GR�����5ߵ��\;V����I�t�?��z����`�9W�5�mw�#,��!;6XTW�{:x�O�˜)�W_.N��Gߺ<Ͽ\���z��'�i���L-�Po����-�e�r��;$���봬��E�T�N=���l\F�m���[�K8& ����C�X=>h�M�<�9l&k���C�e�j��B�B�������p'��5������v2j���M(#��&�U53��W�ݜw���{���#m�N|ں'������jK*���P��f�.��M���юv0���K|�4������[8	X_?
z����<���V�ܰi�f�0����"��*�D`�1�v��\��"�C��}�� � ��-�#���v�7�4���͋F�4��Q�?˗Q%��nw�CM�Ѽ�g�\�p�9Y1�q��ǕY�C3�|��o�薮6�#_ljIy��ts3詰v��E�b'�SH��$�R�����{��ä�5]��Wnv��g��P3�O�S	���:%ԏg��	]ގXs}@���¿-�8���`qUȦ�NXo�vr���;�a$p�B���nX{�P��(rř�����`ӓSq0���4��Kڙ�ц�����H1Pq)t�v+4w�yOf7�<����P�I�֖]��� ��:��Ea���|;��A�(W��eNF�d����|��!0��:ì����l'�
}�>|p>Ku)�,C�����R	1���H���d��<��!e{輑i���o��٣$�����6ƞt�#L�U����Q��&�Q��l3����ρ�� ��fˬ�[���n�e��$.�丐���O!��Ƌ����m������\��עع�S������',�"O'�Z���h���4�	�2�4��}<]hS	į���`ˣIY��/�홟�`�s��$�+-�~3+�;��v���� m��
������L
�����n��=��۞׫�yA��!�)����{��d�t�!�aj4
�}�m��@�" ���j�+�2g�ԮqI`�VcY���WA�������.}�dD���u����>6_����'5F4�|E�s�Q��7Y<ԁv�(��G�f�h��J�.��9|�ڕ������Z#`h�RU% �	���TZ�m�K���1+b��S9��`5�~{�嚸1����h��b��!8�zuB㖙��n�Ц��K��5���$i�/��Ϗa�a���P*\`V��!l3lʈ�=a���}��Mu^���(d�4np�׈�*�v��_�^)%�`f�߃Ì��2���X�KQ|}��r��B��O�~�!4Z��%��}~�3>-zY�!l���H�2�Ѡ�o��s%u�`���g-%8 �|QXlo8T��`��x5N�H��{2?s��L9�� ����%��o���˧��J��	ŗI�)9��D�b�1
BO��,�۬i�{o�IP?.���)g���PK��E������6%J�Z.a��P`oӭN�3\��s�����v�!��Zs�3ʚ~�wl饣�3���`R}�BI�Dx�Y�o!���[�]{E�p�I�č��
����(��q��N�6�K@��X���0C�8\�E����6�O��/ܶ�Z�@ipG⢘)j��2Һ�~��I샆w9�Jk*�xHk.��@��;
 `�p�}��"���6��f�BsG¼��t8�����0��>�bA�����",�`6s�ùXcޞ,��;���͌�]��F"���̾�]V�0�ףt+>���p�!-s'�*�]���<h�BaZ~�$��dl��T�8y�a}ͩ���|��R���m���;�ʞ�7��8���)ƑX�%�I9QjRz~n#���ǧ� ՔtCd�|nD� �5Iq���c�v!"�D�<3���?R�&��W����{O �9�`��m�>�2 ���vۂ�kY�:�W*�;.�$�0l��A-��泞ldNI��%c��ڊb��).=S�Ձ�<g���$Yze��>�?-�~�`:��W+�Q>�c�u�=�nk`'�@���΀��[�(�N��čp��=J4�б����^M�`��G��J"�¸+��B0�D+JD�ޅ��1���y��;����[J_Bd��/�$��x��7���,C׈��'��)�~#g��;p�#�+��mt��j�]��{8IY�Ea]������r�G�)�ZW����+8�U��0�׬��TB1�2F��*,�a�H"�S���h�!~SA������f%ma\�߇�|�AA;�9��+�0���	��S&���	��̿*	@'%|���Y��b6���j���-�=}ܭ�j!���!c7�ª�zM3���w���g��g�#Fww�E~����O�^�TG;F)���-�#��`��@��h�Y�RX:Vޡ.��<��P����yȡ�Ͳ[V}���5?�����&�q�'ik-g�[��]g�G;�c(����O^��S.7��֙?Y0ل��L�=3l�]g?:/������o�FF���ʿ��Spa���9�a��S���i��7�/<��A�"��қ'���z�c�h�XzM�c���Wb�������$�5[�O�A��Ux�~c��G�%�q�Z����)Ps'#�X�3�!!K�����댑�"GY�p-~6:Du*�p�4a]D;8�������m�MG�}�n��	�:�Ϭ�7>@��e0��h���r�n���܃s�}�i2I��� �<3���G��N�����F�C��<��0�V(�ޑ��F�n7^��|�WGZ���'��vY��"�������4�#|ecg�疆E�/�{P�㹫�����1ǅ&Q�.�NN��c9.W��k��P{`m��6�v�+�?�cY;��zU7��õ�k���ǫr�H�/����7 �Ρ�	���
�!��?C�.c�Y��b���y�K]��K��_�CO�X�(�7��X�v��B>�QoE�z�������o�ΨE'���$	�h1�M��3h��{�������K�UxW���}"��K^֭Z��b)Z ��7��ǂ�?�f&1x't��5W&�pL3Dp�n�(�A�������aB�X�Wb�ۋ��>æ�g��(a]��&.F��5S>�y��C��U����j'fpQ�����2�L��;��³b�pZy��j��+� a���z9��S��f$Iv�@L��C�I����`���g�J��-f�ݣ*����������P���z��	-'Q�< 1B�f����D����j����Gx��bű��&~��8"x-ؓ��H���h%��3@K��*���1������o���Y���-��*���8hR})�_���a2Z��A5���l4x�f$���E�����N�쮴a�1��bGd|��� ���+e�Ĥ*0��$LcpXT�yM��=���c�T�y����9��M���C���z��o� �jb	n��A��=4�T� ��D�ש�#P=�w�����XF����Ҽ܈ef��'95��oг�~a(�~���$T*��`��{�2�z;��7�	��o���?�b
ϥ4�÷��y?�>�"�y�.�H���1� ���f+�[�|���K�g�[%;MkT��}�0�b�]��r�
,�����t��S5���ɥ(��RMKM�|�s)�ce������&�}0
����%Q*�*�8�z�6��kB���ٰ݀���<6��fm◑�ML��6��6.�=�8A)��K�=���)rZ�����0�ޖ�&j��P� ��M�i��~APBK��"y�i�+���W��@4����f�J�Weyu2���P�x�u�&��e>?-�9:a��� �����i=fx$l��f@k4������K�?|Ѯy��䬠y?���))]w�oa�:�jB*�����ֽsJR�|ye�.OI�wB7w����i</�_�>XT��|U��:�ۯ�{ZX�P0��������`F�s�u2�(G���/#���˝��?��a��^R�J��w*�����ݘ���U��<�E�I�V�ӊu��!�N=��!c+�L��x��!��zg���
��S�}Õ̠M�9�]Kk>OE�{�<buH6����rW-f��ևF�jW�����Z�[!��it��]H�E�;r aƚ �M�b(hVe��?Y��ũ˲��(�ߘ�[��$������=X�,-m��쭎'Y����ʱ`��*�K�}"��55�q��`�p��8Wf|�:��1U^O��N��5{�Џم��N�D�3CeE+ �RA���O� b�S	���n�?t�1�l���@D�_���D��l����mfğ��=V^��f/�D��=�f|1#�s1�cU�o�k���>g�!�M��HcQn)"���-	q��هO*�T�*x�.��I�ae�b���̋����a�#N��.��ȗJ6i�NtX{�evS1��7q��Xm�c��7�� �����k�A$x��8�ViB�~>�6�,����>������|�D�(���d�IT [ZM޷#B䊟����_Xk'���n�_ӮOq���1�%�I�J��3:UVÖ6���YM�=X@�!Ȑ�P�p���S�ϒ��U�atJ4��*c^ߕ2�5�Y�1��q�Qf�?����׷ S���.�f�@Ej�Δ=�|G*os�8U�덅i���z>1l�+,w��:|��|�/�dO$�r_p��DS:R��R�QΫ�LJE͌�n3�p�*[im�[��j�>4Z,���Y���!a7�����\�(`90�a��U8����eU�]ǡl]�qu�g_�9t�$���7F�W��d	�ǒ�R,�r��k��V�	���������|z&�)~^TK�*(]�-��Ns�(�F5�,�ȕt_��b?��Q����;�-Zn"N�ݭy���Z�#ٿ��E^��?��T��u�!�.����^�����$�b�r������r��wmF�m�&��(��@���#�6��Fɔ9�Rx1W,�b�d|�r�B�ɨq�٬�)%��~�I�,�PY�5��KbxӾn��"���0'f���ی���4�UA�W2sz$C��5�LBJ��!���Q\w1v�g
6B���K>U��4_3¹��N��|N�"̋^ �oԲnxu�+�ec�MuB��eZ�J�i�Wzn�=
�u�Qk�Zv��Qu�y��3Z�)o6����z�X�1�~[�{�Nt�9Th�\5XK.("����ke��S���QE?v����<&�*qVH�vw���e%�9l�%-��V�=E�,**�)�G��`1��vhI����
�	ϋ����y�f#3 ����i!F�א�eZ��+�j�Yj�.Q�f��p�1Oc�T�#���|jv�/)jEZ�i��(n2�a�q�~�`�z��#U#�"�|���ĉ}O���� ؁&)	k�\��M��'F���]�yٝ�� l����H����yK>��N�����=�,�k�����R����`��k>Ņv����\ꎘ^7�'��#j�A�.�J�|F"�!�i�h�&c�u��v�,����
�̯�R�gP| ���C��?��[�*��a0��5�R��Cr�s�?��j���_�T���>������R;��$�Sx�7�=n��5G�\�����p�_��(���U[���Ȇ��'�cux��XY�Қ���& A�Q���I-��QF�=ȏ����͂G֢	`��`�9����L����HE�"��խ���y�*�Y��<�&�b�?��d#)��<0�r�����Bc��P0���lY������E[o�T��%	3;��oC��r#1q	�1RU/���:�/�$L�f���"��0yz�`��]�p-�[�
�u�
`�fp�xnW6y�ўyY&�	��ړ�3a�4ꠗ��d���ɲ� H7�ro�%/�XI.��P�K�+��ᇹ�"�Ǡ��^�� 9_��;QJ��ɍ�&������2���|�,b��-zu���1�H������ 6�̄~���\Xu-���")�CMG}U�-�]6Qx�����r�l˼��,|��!��.��M+/o�I�	�OPߐX�52���>fWQX�%��'�z�4��E�g�0���n���\�;g��A�����5A`(���$�%'�]I��٢$��Z(�M�3�Jo�|	�,�P:�L�)[`(;�ǈZc1Ew��	����"�����	���x�޷�1K��@�w�(�`1�*H�G����;I��*oKP!O%^�q�sFW���xP����Q����6���`�Y� �m�w�c����r�D��� ��%ܻ�Gˑ�Y�!zn�N�4t�T4$t+�}�+1k�{��"�������6cs���Qm�lI�l������ȿl��dKh�K��î�V�'m�'WN�������㙚Y��5@��݀! %�R����(�gE*���B�'k/���̓=I����1�͹�^ۥ�?*�bJ��=Ld�4Hi�Nmh�(U��g��	�!а����/)�#\��{��Z@�b��5�s��U6�u(�a��'v��(������J�J��*Zd�"�\�h@�?cF����m�:�����ܫ���[��1qkY����ҟGw]�@���<wq$�r<5�{C���s,à�I_�@~�Kz~��M��ow�j��`κ�FSe_\�*KUwܱ�bpM+��]3�F�^����¼y@n����b!�����T�i\�]��8t�b��Ac����A�g 6����}�,��z~(���bg��A-x�����o��Ic�9""71���h�3�%�Dp�k�U����G�h,14+� O|X�3�o�b�����-���Lw^��\�k�Zl�{h��ԕ�@��u�I��A9�k��]��~8��z� ��UV㝜mL�մ��=�Ã��pR�Ǡ�@��4�o���<�r�N��P��W�;�,�Z*%b��y��o��[2�,��xH�T����߭�C
㜸�8l������뺾��?���q�<����la�6}܂�#�Rs�BU�^���a�j&��������unC�QwG��3x���ɪ�w�D���R��`�t$T�B>�2de����jÎ`fN�`
E�)O�	R-S|�����$�P��	M4Β�	��5o��0�;	t���P��$�M����lR���/�dO�O��9��dyx�W�,z��4Ý�3*h\	mG�4EU��/o��<����&�a��*L�0�A:E`�h4������7tX!\fAs�9�<o�Y����!,YE��:({\�� �^ �5Y1e��P��A.S~����毥�OϿ�]�σ$���O���YQ[����A�]��w�������Ԗ����8���n��E���F�!��+~�	z��]���ߧ���D�R8jL
���`K.)�v �Њ��a�~��!c���̕I������z:L�#\1܄/�7�:j���׵�>�θ�TЅ��/N�m�(8�d�Z�<({�����<Ni`�)X���
7���׍�c[�%�d�T��Đ��1tɺ5m9 �09�����J���L�nÜ�U]�,P�j�c�AE���zp�԰�Q�Z{'���� �"���R�9���`��"����|�!^0�����F�!��c=��{���#9�֜0��cc��D��;d51�Ŝ�e�5����[�v�!���pbGbw,�_�$�[�qW��NSč�̾2�9�1�Ѡ'�ߨ�o��O�k���s-^�>�C��ئ �i�+�޸��P%�;q�U����>#���j Q�e�8#�m�#)����*�YA��L���8��j�.(��.T!^G�Xv:�s�`���K`�L���- �}��0G�b�V�����A��qaB5�@���˾s���G1 s�/��k�f6�+�C-��3�9wI�bH�ntY(�:�憹��s�4�H�_3������Kk�t��g7bɪ+�z��}�5d@	ۅ�U�z	)�E`'\���_33����H���u��$@LpZ�X|OO���%x8[B����bܐ��R�F�9"�J�����;&���}��G��p[D%�B}%�����T�<��[�|�Y����0�N�!+Z�i�~���A1�u��<ȗ�Y�#!�������He{3)���Pq���_P����_Y�����>�)i'R#tIP�̻�,��ۣ��ONFW���ě�6���_9!���b�Y!��U�j��y��#���0P�<�~�|��5?�~Q�����Ѡ|��7�z<�'P -A�Nt/�_b���*��jC��׾�#�5�Gku��>ͥo��՞Q#Zr����c$������ۖS'j�Ê|��dT�-Uv�Mƕ��!D���+v����E��Q�Q�^kG�0��1O->t�PMϚN\��py�~�h��cݥ*�13�?���`���,���R����=v����(a-[T�MQ��s�$�0����Z=_OE� X�]�w�ō|Q���f�]�|���އ��Pa�G���\焩=�*���Kr��O��7�b��)[�C��X�uh��	����`���@s�W��O�w+eL�Rp�H�^3c�X��P6��r�%����\�d���:��5�Ws��R*�_52:O��
��.��dd
�`��W~~��قl�ſpʬEl�U��?���/uUS�14&��4�������|�C�&��a�C&��J�i��k%�y���\��A�'l{0v�dԉ�V� rjK�'	�*�]��?�1����Q{�5�%���!�h�^Q�$�9C1�#��N���!�n;^l��]!�E�P�o�eGq�P��+� ��ߢG����FF˳�b|W>�:=qs	}�&�O�G��pJ��yi0�����0y���������{�ԃV�#`�����s����l"l�M��2| �K��������qf��f(���b�#��b�������2_���S�v��u'c�k�����%� �h����ˉ�Wv�O`���GW�	L���W�uf�9�v�vR�Z.g@�c���Y��	�*.)���w�J��X���
��m����j���T�?6�鹶3��"��{�?UD�P��#j�Cn_d������m4T�l��i��,�X�I��:���G�Gf�9�͛�z��R�V_�� aH]X��kL;��4�;L��hYӖ��|��bb�L����M1c���fѕ��"��ܱS�����(	��u���3D6���(A);Y> ۋ�r�&#k���ڿ�L�݇��*>��(	��b�)�5�"��Y�� 7uȥ1i�i�3�X3�;���*4���dgC"D�0:e��l���^��l���dΆYS�#�ی@���h��Hs���S��j���.@Rq�-#�.�eb)�m�E����H(CS�����H��M&4g_�-J!dm[��K���p�6���?�#m{J��:�𢞭�_�����v��Up�9���m���s.޻�t�h;@V����.�R��#�����0ȏ.��*�.kH�;~��H�M��nߡ���mJ#�¸��-���s)'��
�TG,d���pKy%BE�b�>s�t�R�<��hQ#�=����S~33u*�����������v�-�Qa-(������j|��x�R� �@H�cs�\�P�ϓ�@%f����sM{�Ԥ�3s	���ra�[�t>�娕Q��N���u�H�Ok����?�R\ˡ~�o�I���3�"��}"��ږ솣7���5��B��)��àʅ[��)Bʞ�����)C�����?3@X��)"���
du�z����R%��$�1o�/|$6��0�o���]v��"7��$�L���6��j�:H��$���4��;t�j9�U_�[�Ψ]Zb,R�~{k>̯�w[�^�H#���p�d[��zr^`y�����D�z���@r�� �LWz)�A�k�e3�ь�a��������Ͼ���c_����[Ʊ e�i�$���u��.P������͏ywy6���2�|S�� �M�G�Pi�u�5Ǵ�~;�R���ʯu���I3�$�B̕u����桑�ØZp�H�YM�-s�1�-��g�����J�IE/́Զ4�{[�O#�HW{��SN�3��c���Ƞ�M�:ϿI�z�`��l���?�]xo��r�ř��~<ΈJ�^�z��/�H��j&�5��8���7�I<mh8��Ӌ���
F�֏����ea�t�V��x���{��tY��dT_�7�7QF�f⬰�_��]�4Y�.�����"[)M^:;�� �S[�w�j���ö�j�`������ge�wU���6���t�����.�� S����'��;��v��8H�� ����b�̲'�8�2�� =�h���~�J��VY.bFF���M�({�ƃP ���&�B�nQ�_'��)���EA�~'z����<А�H����z�aAV鿬���8N�7��`i�-2�#��>m�`�a酎"�(��U<w1P��GM{ �zN���5a�٥�?��̉�X�q�T/	 �տW�:�~���4'xFse���K��)4�G�j� N���`����k.�u���sn���������к�$��ϴвv4���OJ*�b��nWr��U�~�����Μ�ɦ,R߭S����a��|J�4畆�:>!�gh&�%��(��Hx�GR�Z4�����k�q��ڙ܏�'Fl ��&w͌tx�7bT�������+Z�;M�W&�9�R���A�~���$�*�笓z�M{�bQ����h} ������w&�d1����$G���V28��C�({����5b+U�&��[�{n�p12�s@�a-�
��I��CF1]�a���Q�׌�}�a��:����3�~�K���n�J~�G;�T��l�;%�Gxm�T�> 
�x����#ԆT@��/fh�>�u�"���k6�U�<��i�-wLyz{'��v$尦d�����$�C��v������	Q_s��'��1�R���$��>���Ґ�+����!��'p�V�BP��P�����ۓO��?}�Չ�&����d��Y|U����g�?���V�&���Yd�R�xg(�Hd�!� P|�v��%�߽"P�O��V
�gCڵ�J�:#�Ii��փa�P���(i��\s?�`�0�@4��z�F����x�Q��c� �?x��3�n�H��|�g�|$����������z����>��w$(�n�Y�^9�8��}���ˀ�!�������5���c��%c�6����P��}kt�*R�]�)یl�*YhA�_Ȁ#!ޅ��G�ҫ���y/�6�+�>[���:eXn�<��$���m�/2�]���A���6!xr�J��x�8��˄o�y}.7L�����q�� "w]�<w,M/��0�!��2o�^���ݔkO��~���IE��c_o��ٕ �,4�k�a��Ð���u8Jj�,���ۧ�b���ڛA�l��xæA���5�֘$�Oj3d9���]p�./�
]h�6�Nk�'+�Dn�e��|��	�w�l���4��WH���{���;	=0�N21�4�#�����l�hү~W��U�W�?9q�zd3����� `�D/-co��hP��.X�j�����sW�P/ Fo��P����|����-3*J��7E��t8-1���pq���i	.\�R-�E=;����o �A�{eT��Z�=�:R���:L�:�R�b�ϲpr�ؽ[���\�7��KT+Y-gϾ�n��l���~.�ofI��@�7�IKAk�8�d�����Q/��3Q�I�mn��=�Y;D�UK֚�ݱ��M!~�s?N�A"Vgj!���-U��k��MMP_��?��f/!C�h��c�}��V���Cz?ҥ� (�3��Xk�q�|�ȋT�f����\<��zё��V+_wT
��y]M(�������K�����F��=4�N|K&}�u	�4�vHA�`r4�̋��p�a�6�@!� P[�AM��S��� �p���d��k�����٠i���w��L�8ވ~j�PfRMT#��5jt�2j�*;RN�ŀoߩ(��+�k�Y閔���u� �Xp���r��e=G��4�p3�����چ���&��8�&���\X�q�����T?���m���)����(DK�KL��&��ܫ�^U�r�D$��A.g����j!I57�:��'��C:��.��o��|d�����5[r����8(R	@�>�j3 ?����ˢ0�����ߛ�3瀭���#����nDa�ܣ�I��6��� w���hP&���v"�啮Ũ����]�|Q
�1!��O��_JX�/�w^XtBP�C�����$|��&���Pb�I k�Wi샙�-<���Z����%���_f�u���QA�|��<ЬH6�⌛���=UВs��s��{\�(86kX�2+ڹ�m�$-Oe�\�K� %7�5"��VӣќT��)�F������������:#XX$%��s�(�!_��]/��d�����b�O��g��x��S!�(���vHʀ���E�W@>�@I��ɓ-���Y��z����(�V�`mm[�@+��lNmct�/8��0ɯ6��.1r��*e���%:?*������
�=PIU�mKy#�������xx�d�УI�t����7�÷��6�NC��"�$F����^������h�ТHidu��E�F2�H'��k�/�]���p��9�k%4z@"���1T��tr�-���>������1�hE���]���KX)��6ut�JI2�6�nmWh�F��I��Xd$�J��\(�(�c��2��j���A<~5�b�Î�,1��+��)���G�"�?�8|��?��zyFl�O��"�u�e����^�#������P0�Kuv��q
�|LĄ�j�A�����ڽ^Ʀ���@�M�%�S=ۣ�~�'|36X��)����Ȏk�Iut?	$�d�k��(t�p�鞶�������;�.�B?bg� _LV��=�"�W��R6��%0�c�/���l�iَʞ>f��R����9݈A�K�<Z@�/YU�a?Ar4�,W��q��
�S���y�#`�[� ��!@��f�{�ƿPG��H`� �?>�[$��/~�K�!�I��%k��[ܕ��?�^x#��Cs��ec%�s*]j�*A]w"�O�_��iy�ӟA͡FN�x��E��*3=��R:��.�A�*M�y,tv��Ý���0f_���<�S{����X�^pVlmDߑyD_ʶ1���������j��K|-��#��<F{ꂁ�����5w\�ۙ����g�A��=v[؄5�dfY*T�>
j,o�U���aq_vy�C���	X��^}����g��d�c���.\~����5bId>.�c�z�}h��?c�����o�+��-�MN ����o6���T�S������B���{�����/m��Boǳ~[9�����N4�*��ˉ$���U����;��n�O���1�_I�h����a[b�Y{K�C��g$�3��$��%���y_Go��sn��P�kA>P5-f0EcԨ3��^�u~bq�T�+č0�l���|����c`'�Ǘg������|>#���l����ه�e7Ǝq�'�4��������"�q��`�1�����Z<��AB���~8��� �[˃����5�I[X�'̨q�y�Z�K�벹�8�- @�F\ǳp�I��׾�u��wM:�l� U�_Ay���/6��"է���6Db)kq����4癮��0���BFׅ0h7�.csM:&kU/4�8I��ϻ_=�?�!��Ǹ�Rp]ˮQ�WO���}�0��'Ǡ��E%?{w����"�y�yk%F�f^U*T��y���t�߬Ҥg�3�8��Jc7�_Ӡ|M���o
_E�b�,�G�{�ef@fQ�9���b�c��y�d$�{yM��6�P��(H[�P�ЈnK����'�U���S�d���?����5$�o��tԠy����V���\X���0q�-W�E��,�^k�p/�;�-t�p/`*����p���rC�;j�w	bS���Wv�?v:�ր�d4aW/�ƹ(Q�#��5w"�q��w6V0
]l�b��r�.�:�/���#u��<J�E'_[�#ˬ�j� �C�.4�#���F3� v�I%Eo���Q:5��gz}Z6F��â�r$�7�5�k9Yb�j�>��>��q����2�b*�Fx�\v�ZRZ�������:�8�6F�qN�<�+��c����jQ#Is#�'�� ��lƶ{rL�_�=��[98�j-�|ɡa�Δ��^��s��֔SՑ�����ePa�.�M���!�c��ٓ�GX�����BM�?�y`5c��7,я�XS�D�׌O8"�ǻ�/�8������Ju˪��Oٗ���'0ȑ��,̪Hvv�A�1H~'+8l���P#WwT���ݣ#���B�w��ʽ4]�p�Ò�^���j]������)u��0�Bil�$�٢��ڿ��!��=�;�̆��ز2�����Ջ���Y�I=4t�����c�Ů���O8��	� ��s>�mUwAz�SMi���8gIJ�L����E��"~{�_q�e#�G���G+M�,a+rl���!������Q+�S�j�-B��ux��|2�r~��6!�[��UWx��L�}�Z�1-5+o����X@��8��ovGÏ��0n�K"s�����r��8NvM8w�#�Z`��O�������h�pq��$W�+FM+ 姟�ְ��-�/�t� _J|���9ߘT��b�Iw� M�"��9���+H��3�M�w���J֘�=*�=���E�3�����ĸ�V���Ͳ��/ J�a�)�Z��@Ř�W	�^���LoxvSֵ�~Y�q"�kyS[*�DH���p�]]�`�4پ"�X�� #�2ȇ���d&ܛ+G`��Ď���O%�Ȱ�!�!�#>�A�v7IEI����ܥ���g�cj�SZ�ɪ<���L9)�EAH/(hS�[��tLHs�AhX�3��.B���S}=z�v���p�l���G'5�]Ku0n�<�t%��f
�A3���8u�B������K�?u�X�@
tq�R�^J�`��a��T�٥�f�ڢ�9�߹PX0S�GD��
^�'e�����c������}�Ad�V֕��b�Z�����rGk����t(o��.ΥaϾ2���[0�g$���2�"q�V�HV�9{0�`�5檎��{ �z8`>��+�o����N	U2
;�i
�C�N���]��%�YޱYO����~w� ��$ԉ�#�в(���k�ԅ��]I�['+A�>Dϱk�A���{�wN��/�:���|, ��W��(��=�C��#1m������!?~4���-�v���?[ۛ���U:�:��O+�\�oO����5��ۭ�N(Icrϕ����� �,�k�Ǥ1D��?n
�g ���O��8<�� �3�~�.J�mr�Id��	�q���Q� ��E`@����Pf�$��^̟&c"�l��Vz#C�l��n#�����t��ҹ�aP����@][b�$�|avAhA�Os׷��e�� ݇�@�W�F$�_��N�gK`:0N�Y��?|Ռ2�Y���DQ(���Q�k@�qC�xZ�p��%�3Ϙ�!�t/�Dw�D�(mA�y�� ����yق�i�:~}�9�r������Jpߥ:z>���A�y w��3��pN������d��G��*���JV� ?+,ITp�]ǥ�
�_z�>��|�|�e��wb��f�5ޣ�t&�2!�g&�E�:HjcQ`U�JZ��m_6$�� ���(؋Z:-Ix�� �O�7?R?�E�!G*G��u~����-)~�����NeS<��v�I�3��N�1t�'fi�`�# }�wXÖ-q��,�*"{����������� ��!��R���P�5ԭ_m��#�\{wn5��!-�"�Q,G��y����(̷��tZ�i ԟ�S����&O�8/�j��� b?�۶��%Qu}�U"HX��[-P�օeֱ�Ǎ�{S�ݙ�'�G�w@�Z�Ik��P����Y8�vfw`߾�� ��d��;��r�x�5v�Y��;Ц)Y����m0����r�Ǥ��J����My�4Rҙ�wM�")�9�p��s%�� w3a�5D�[%Ԯ�dX@�K��t��S��n&�V���t�C@g ���k�t�he�"��I��ǁַ�W�(�i%�:�m���žX�#���"��xL��d��ϋ��/
"��BQ�Sh�Sp!h�#��s��.f��I�OM�踸�{�Ό�Z��X�A;���=�����^��lfL��]��n�,e@�(vXteUPR^ 1����y:XCߦ�=�K8,%�Ø�m�O�7�m��R�f�ՙ�؉%X&wu���a��2S@y(!$^s����}.�\�y���d"P��<<XՖ,�����>P��NӸ(2��JA�-a�e���9A�D��jfC�'��b�u�$�g�]��:��D����>�S�^᩻��;��1��6=��Zl�U+�pT[��%$>k>�y��t9�5�~K�9H}H��[G���;�W+͡�?}0f��Ϭ���8��c` ��uv����u�A�&�3��n�;��@A���ǷI	��Z����g�W���%�oM#T�5t����&�<s�(���F���i堓?ѓ�ǩ�y-C����ܑ���2�Mk
K%Bk�m��y���{�FYF��~Ky�W+�u�r�-��K�h<c��B�L��5�%__��Ua"k��jpV\�J:Z�iq֏��� �ʠ�ψ��Hv�P�Ҍ������a���†ȹ6p{�����F��k�Q�\�
�`�m�[��U�$�����]�^9@�t%�n�k�:����,�yy�y�,�oB:5M�������3��]�-�G�Ƣ�l{�ݗx��z���Ʋ^���������b���^?V�Z����w'��.@�Zp|��-,z���� �B��[$'1Q&��$=:�N������J��W>����ZQ������4/к����B��3�x+�K�s�`����E\F���@�,O��tpj��,�ﳉj]�]�A;�7�ń0��6�	1�aX����߄e��>�pLX�y���6ܒ�妉8H�'��{2�N��;�<�wq2��e�&�u�^���Kڊ����̱�r{�YĄ��a�$�1��i{bz�v p����U�2��z(fWڊ}�!Y2��(�?	��Y��L��{FXC��9����w���4��߶�^���sɧvד�G�(Ki�,i;H��h�e@&����@>K���z ?�����IO�e�o��4�1p��'�oK��}��xJ ��*b���:6!h�	���@rZM���U0)q������j��T�J��w�_ј(1T7�L����ϳZ6�=��5�W�7�s}7�k���5�FNj�^�|J�ѭ/I�!	�̬�AeI�R��|jQ��8YOpRK'�]x��#J��\u�3�6��d �f������)��=�9�;J+����L�F��ŷE��Ů�����UDP�I`YdAHՔؿ��%H�!0c�D#Ⱥ�<qp P6 ]���7�LB�g��'j�z�D��^�.���
T8ǗF�<��|&4�h��J�"��g�a% ���?��I��#h�N�����QK�%���$I�ڑD�����yJ�o����3BN�&����1ht�%Bw,�óՠ�x۹�u��yS�XN��F��0��-�F�v>����̘�	p;ʗ�^{�m�~/<y�F'7v���'H�ٗ�+�l;vא>� і1�y�)<�whi�wuE��ٽ�� �ܦ�Xn&l[�͓LJl�{X���}_%��ܯ���Q͈��Q����GrQk�L);bԟ*��� N�C�G�������d�|K{h�R��r�x�,��Ȳ8ܘo��#�5�D�}��R��5
���?�m��)q(M$Mg����tH�ԥ���s����7z�֩/x�Ӥ�X�۷	��82��Ա��+���V-�)�X�3C�]�j����W;V�zÓ��p�o�Eu[Ī8�O��T���3���b�=u>��7(p�!pWc���#PƥN�ƺ�lȗ
(��)4}ѻ=����XV9+ʩp]Aq��&F�4�'&�l�;,4Ԋ���l��zdK�[��#�E���b&��Y� �X�]q�ܾģ��R����a�UVT@%�(W:D�wG�nm`�z5�bయ����24��sCÏ��X�z̾�rXvBIA���wL���v�G��npI���MF'}��t���Q��X�CP���