��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<��]�55^4��ԇPD@�?����Y�ͱeɪ�N�uQ�l�>�F�҃�R�yk�x.-�jeCQJ��kXY�os�Ca�f�|��F2�Mo�4f:������H;ȟ��W��q+�,d^<���	���(A���J��(]�?�ҕ�Ѵ��x�b��s~i��:rQy9���[l�)��W����,v��?�4AW�v��x�<I���'�[(�=����_��_�AYH��'[-�2P8�)�։|�F�����u����7��"�pU�%Y�y}�N��mjz�	$�(�"�k/�,m�Mr���G�ӸI��B���Q�@�
�÷� b�,u �UD���0�I�`���H�.���C�.�����C��&k۴�JvzG������;4����~�N���J ��B&pm�^p�K!BKiU�ab�!�O<|�������-#��P>�M��(3���r�ڵ'�x�
�����_\�k_��Ȅ��;!�΁�6�NXPhdm�kky%�#�h�W��4���H���|� ?��=�-�+��^y�"4}�tm�ˡ�k���a�T�'`��l)ICC��,�k4̻���-X��uC!�����z�݁}0��s���.���Q���	�tk�3EbN�8­�`�l����p`K��)�(;��p�<��G�e0������BLO��n����u�������C�;�������HfO��&�	���b�3�H?�ﾧ�f�]��.�|��#���T�����j2͹�)q��n�6ͭ��z��$�[�N/x��-�Hi-�_'�FR>g�ZE�`\��J� �D�HY�up�D�ht��m��Z�h+(��[u%�����]�~E�MV��&|U��R� r�I�x���|��F���w*09���/��j��ע���c�{�ɲ���}?���/�Td�_E��^u^/W �6�/q���C�Bs�?x1��ԛ�'^>��n�q�թ�4���4Sܮ��N1��'�on�,���%�5~�Q�S(�������q�0��p���\�#���3�7���7F�8�	5�#���2~��w�p�;"�����H;�&�J�*)B:�F�s�h>�©��_j���-��b���G���,a�%$݄�Un�nk����|����gߡX(�e�M��	^V����u�F���%^�,�X�a���J������4�V���$��cCբ�fAzdp��noK��1��J��|�����a@���ё�G�3%_=I�G�K����'b�����U�C`/�Y� �P;����.'�x�٬4�n+Y߰���5���u����jx�TzZB���E�{m��ԟ���J�(o2w� ��M�Ƅy�+�}� p��?E������)!fz�"L0���cd`N��J�n��0���'�z�r��T]����a������O�l.;�8a��U�g��0F���뎘X��lQ����C���[&>w���E^�<Mg���~\�2��.
0���.Yb�/T��=���؎&�D��m�C;�%�QM6�R��kjj�9M��@��@
�z',�h��۹��6-�࠱����_&Ӡ���a����B6�8���%�� l���驌$`�K��������>��/�މ������~���6�V���E������j�`�ђ!S�
���p̢�7@Q�y��ޔd5g�r ���I����n���=&�����7�2��-Wq��SӯZ"s�!+�f�<���W �4+�T�+ �!���׮��R�]���TD���-O���{&ۃs��k��}Da��5�̒�D+U�P0WO�]�|���W�J+�"<�r��fhY���O��H����sF�Dr��R� SuZ�w��>I1���M�^\��O�!BM5���+��@f6�P1���\��虊��]Jڙx2�(dRM�~G9^�"�eW�`>ޣ�ѹ�؁6�Q�A�A����bI��y|mV��3�FJ	�ᐫs��E��Z�d~��-�ǥ�zC-�jzW����@f-�	}�⤸eɺX;��0��	�>]GT�-<�eL?�{�f��9������M� ��F/��6��
B7��2��	�=n�K�jR��WV�����N*!��K����a�#M���|�h쒿��!*���Z���`��+6X�v"Z`�_�<Y=���%V�_y;*�F��gX�V��s ��n�-�v�?�#s�fG���7���F�ڱ���M�۰F^�����&K�l�{���P�=�@����{F��W��Z�%r�-�mN�O��=d�F�*Ĝ%�F��u���"�G\��%Lk�!�'�� (`˚��!1����0 ��P��-����?iI�ץ�Q��XbH4����Pk�W�ɳ��^��3�X���0��nw���'=J�ӧj*F�������7YA��|Gw�h�ɝzJٶ+��������ZZ�Lȭ�F-���0����f�7��