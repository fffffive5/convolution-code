��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L����ʩv�*z}	�8p�^l_+�l-+ӐǷ*���dp(<�+�Xd�J�mT��ga&O���C-�����k���.
W㓆�����<�Z��*Oߜ���eo3���	4�K{��,ez�.T��e�ke/n��\�����������h�����<s��i�j�Y�!f�}K��MȪ�3z{���<�rx�t3�G'����}j\�%�������_(�  ���
;��]L)P�ki����3���j�C�,���N`V��v�&���'y�i�� ��[漯�S�0̌e���h`KQ�yjdLϗ�Be�;3��pz/}He|[{9�u��-�����'v,35���q/8��m~�B))OM�!��8����j�\�N
O��fr��ˉ�z�Gq���p�3~K���C��.|П�J�VlX.4s��/�?Ú�C�&	���T�#�]�R�7�)�@O"L챃��� u�f����C����D�EJ��.m����C��K�ɮ��qQc�"-❹M�e�(�w���i< �c�"*\��-z�}����w3=S>�nlh�͓��ܳR���|}�L8�*IK��*Ȳ?Ho�]�V�򥊛��E���p%�vy%��e�9���*F�T	����sw
LXB�^�/i�d���E/�e��2ќ��l�80_0��s/5���Yi��|8i�������@�]f1��+կQV�t�yeS�����������T_�˘A�����^&T�Yp�}��rRF�*5LV��E� �h)Q{!�|�����ܲ�ʙ��Hi(�D����]�d_ZB%%�f�1ƥԉ�P�>�8�r<5)|���p\�lz_MԺ��������f��D_�����Hv�4�#rA���?R��'��|>�a& IV��u>MW�U+K��xo��]��S��gĮ�j_y�Mc�-��B��`��Y彙�|'?ybV) ��H�<j�t�Bg21|��Ozx?�"_���� �i�>���j�pni�R�<�β@�K(c�I/����s�G�T|�ֹ�y@���4M%^�S�&��������5���g���C^8�]eȉ�+E���_�|z���ү]��oC��%�mr�eӂ�Y�<�+n��ɬ� }У���)�Z�i�z]d!�?P��� �
&��Ih�wk�)!�!B�ߒ#���L����`��5�2��q�-��/�&�ҡH棭$xlxV����g�ҝ&�6Y�s���G���D	�;n|��e�m+	���{�u]c��Z�&���	�	�\�a�Bg�,�%u�������d��n�c���%{O摷
��t�įa �%`n �\�A&�;�ihRB���*�!���7���g�8	��#�s�j�� �1n.�_Cw}b)d����Z�� x�>�T�H���8�6���$U��M2o�#� /��:^��bU`�= ��@]�Br�`ur!���=��r�i��k�%N�y�����#�8W`�\�Mf���5��aTv��Di��E���