��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<��}plS��w�(E	p���Hn!M�����!~Q�Ѷ��0�+���z�f�Cp�U�G�x� ��|;�������@����ܗ9[5�V�H;a�,��nv%���K~UO!�uiE� p5�؆����L��5@a��ڴ� �c��/H� B�gnM�ͦ�9�
$MW�fi>T�vc�q-0���¿}�L�E�4�SE�EZ�Z!D��_xyl?:Fվq<�G+NͬE]��I8Ҿ]��t~�h2�v������Oպ+��0�*�.���w%���3)k�S,�"��7Ix���0���I-
6�Z+����4D�ͷϮ
Z�l��4�ߣ�<���c�+�I�>#�ұ�m�L��Jݠ�Z5�����2�'f�������n�g�����T,е��mi;}�4�&�M����Ş~?!ڂ�HIi�x��>u���%�$Q3ʎ�Ċ��/p`ܜ��3��q"�ws�g��̈́��}b]��ɲ����n;K��p��q�{�*_Fޮ�`�̢�6�o P�;�e�����9�.yw�,��J�~,�Nmlr�z٨��
Q�NQ9�y�hXd�N��_�/ ��n�ۚP`Mf�N�:~&]�#����D�U�Ͽ��������:���lP��ǂo���E�����Z�T�_|��U~��B���W��� �u6B�;]f-.S���0I3��嚛h�s�ӓŅ��b�|Z§�� ��8���
�E��<���{�����(T�r�1s, s��ґ�ֽ`E&/X/�#h�	O�'��A��jc(-����e���d&���G����6Y��I]pf3��]�F�d5ήx�<hR$Y���E���6�b��خ�F�O*,�����r+�\�HA~�<d-��&����g�����4��{I��S��`��Q7-u��h.�'&�Ei5@����o����xTNU�I��K$HZ������FC �+��� �D�X�##��~��W ^�<w	��pao��)�~�n�_�W5����w��F����3�yy�i�n��h��/ӓK��($q�d� E�#bt
���s��ve9wC߶WM�Ȗ���8�;����M#Q ��Hx?��H����CI���X�b��1���������};�(�6� O�p�7k��/��G:;����cuv�x叽`Й���_,�ٯ�4_�*��<��~+���ͷ���������z�������V^�2�A�Z��;E�%0lL�"Aܤ:����������d"���{��n���qq!�hC�v�;�w��961z��FԢ��}��Ow�q��	f��ת&�a����~~��z�r��<0T�?������P���yJ�~�X%�.�gi��!?�{̂��F간{�"d|��@���K���s�$Ϛ{n��k�=RH,HW�-HE�Cƺ�1��%+�����f`'H`C�3K������/���O�S�����룣��MX"G0�R�Ń�)�٨���l������8�Q,iT�n���jh���
�١�+���R��#tCk�����@y�B��-Q�q���>`"N"`T�!N9(�EL������!����NS��ǎ���w�2�@��]){F����S�eӃ?$i��9�%n�����v�����~Y�x�U