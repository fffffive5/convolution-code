��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L��w.�g@]7o�V[/��)	r�٨����s�s���"5����pUK�D�����k03�e~�C_u�T]<��hs@�|��ٛ\�1��!��E���w>c��F���I�Vu�Wj(r�Z]9��:�+��j�c�#��X��e����̖�щ�ݓ�z]�����~�B6�P2x��&b���,SN�������U�T�C��t��,	�hAq����"��� 3!�䚀���($g�랍c��q�r�����¾,_�,�x+�mrdi��;'���:���pK������ή�௭pq����g �wD}ɝ1�c����"z}��!�ZnN���N��;���ݦ~�O:�q0*��J��ã0ב�$�6:P�ģ11��#+��$�}I��\����-.d���h>���?�x�h2O"i��F��uM��6 =(bY�tk���u6��#LB���`����qY���*����R��!���2�ke��LK�{Tq�݇��œR�͕��¸c�/��q-���+%�5�l�+p�R��P��"��c����Ԅk��?Ub�VtW����;
X��YՐ+Q�e/4nw�P�
�qbYߘ6�SFu%h���M-�fI�6��L����pHs�t��I��5�#[��P�����!R�ڙV���b��܋Q�*\z���%�4
�x�">��J��D x��!IFY+x �9��Y-�-�?n5_^7�Ǽ&aw+s����86J��C��-5R�؄�� �Y� {�����l>�����g�ײ�gg5D\���>���Ïq
v��?u���NvOԺ��*�����?Ȧ�4l�>{��t}���X�� �ɷXZ?�2|�6��ʘ��`o�j�1ܭN�2�DdX5#��9��H�Q�o�0������i��	^�V���i0�y��S�}yr�$�&��	B�+嘤�k�����ϯL?��&���;A�g �`���O}3]��uPY�9'�C���w�٣P��8�ҫ�Wf~-�hL�*S͡�%�6|����Ā����A�'���4��p�v�w��FMm!�--�+|�7��5a2�|����N.��,)�p���b��ƌ�����96*��Z��H�+CS�{�w�<�;��i��7�S|�Xۗ6u�_�H[����A S�S���j^���x��7Q�f���_��hGD�=�ֵ���{�ݎ�oov-VF0Bu�g\=�o�z&P�V��������X��"����Sǯ�7t���e�dʱ���jۖiB�
�އv�d�K��\9�^j��<�	�=W��j0�3I���I�3��Α�B ���������9���<	K���������Z�?�-�� ��40�Ov'��y�w�䠭���{cE�*qv���힇��A�m�6��k!�!�Q&j�V9�� �M��z�oX�C�HfW`�n�ˆyq������]>W��j����-�V3HOe�T<k2�h���v�@����T�?X�����-��#�1�S�)�����X��fMC&��{z����M�)�(��:��S�Ju�'����.b�� ��D���#�az+��z�a>�c)�D7�mS��'P�Z�Y�K�Q~vP�	������q��k����"J#���.��}����N6��+g�NƂI��w0Rnͥu���)��C�O��%��E O�S��#���؊�ݤ�!�J(�t�x}|BPvi8���p,)a��,������7�~VS���>\�3FSs	rl�lxe <�mm^���%��5���g韍�ڽ�3��_y@�ղ���`�2�C��_�f�
Z��f[����3���utРVp�Ï��j����pzdf�f�@P��
�o~a�Rwb����}�뿗�y3�-���d�z��VT�^�a�_ΗBl_%��*�k�[�'�w�%X�
]/X��@O��X���X�Ho�E>���N`_Z�����?lx����b��)�a����3d�9|����A�ȥ��D���M�#��G\�F�V>�l������$4����ʆ#�y�}_��;�F� �����m,��qb���W�qvno.S��Կ�mL�.�����87��<�{=��X:�[�gHsXh��iP7$�z�&�*���W�g]�Y�3O��QR4+1��rL�(Y�QR�o��ќ�7�J���d��M��CI�N}`���L;���o�)�.��&�]p|�蘍%����Zy]QM_�Z���a���K�50�PM8W�����~#�&�������d] 9����uM1��3k����·S�Xȁm��:x�v �|�9ݙ���U��Q��e��`���J�,�\X^�s�Ԉ��j�Չ)�5M�vi��@�i?��f��lܹ�I@uO������k�k$@Lg���(|W@5u��+|A��?����-�.|Ӄ7ܻ
A���T��B��Q��G�ٵ��gUV�+�7XT,a�W���E��L��x�iڪ�P���d��A'��
eL4�;S�z��%�r�V�MCs��=
	���Ֆ�E���+��=���*n�oJ9�����Ԃ��[6�ʦ$#K�
l�:S�Xflx�I��t~�`I��ѕ=v���OwJW���N2i��*6�hC��"9ceT��D?Ŀ��L�
_���s$]C��_8��Y<-��\釜$�;�ǯֽ]�0�2���Q^8���%�U�z�}'�%��r�P=��b���q��5���^;���u+�>E0�+��Xצl���Z�>"�R؀칒�/s��m�3u�#�$�Xy��a��qc�5m>�?���4�#��\)Z�JC�5���S2�nN(�������@���+~�� $!^UM.j֌0�!~��y���m�/��z�R"��ƤH�`�x�Z/�N]�V�\DJl�S���w��z�]L�ҲQ1W���:�:<2& �?[�5��)����U�M�N�:��c�u���u)��F(�ʑ	����Ui�}y��X�22j �j�F�(/�֤�>�G��T,��MF4��J<��PQC��/Ϛ�+��^��i�v����I�Z8�$���d0Q�6�[�����p���y7ʬW'���	�_��(`�Sؚuǝ���t�'c%%�4���]dg���ekb�G������I��;��ī�@�͑m�Zjv���؂�x�sCfE��0���w��5]_r"�^\��'��>���2N2�����ktWrRf$OR|�t�푛Y[�Π�"�ѳ�D&��Z"�Q!s3���Ŷ�+l�e��J	K8�G��M�f�PUh�q�Н��=Bq&۶ʹ���1�ԧC����4��W��,���ŀ�+�A��X���{�k�׻��C@�_ӚE�ϻx�#w4 �+REї���<8�K&�e8��^�I��ّ��6N�o����	Ҥ��.9H={�������2 �p�D�Q���5]�$�d%N�am�6����>* �Ml2������Xf�a��tRS�{r�M+׍W�P����h�%�_��Z䋡�d��W��� ��G�y�7��%�x�N�ՊɆ�C��)���^>�l�.ݒ�{�5���7
��֑�o��R'��|�<U�W8����Vr��A�&���Na�L1+���T\EQ��^�?s��W �V�r���i����?[WR��M~.�H�g߿v3� i��"��ɒ� �Jeyd��v	�"O�!��z{�>�э
>��f�3^z���6��q�Y��*��;�p��8R�!o��gf���bF����f�2K��n�)��[�3���Ȝ���$�E4uY�*�gGչ�s����5�{ş�7m� �I_G~�t��i�( �Sc�aS��=�b��*.�54s@���V�ݖ��a��P }9���a}V��	!�O�`���%�-�.��=���t���T�5nX�Bw����"c����Ք3،�'��H{o1�1x�ʼ#�U��b]Ӈ�oGl��BPٿe�,^�D�`�\Il<\b����0� �L�VSߢ�̋���aZ�x�SU��mFY�I��7PnZ�� pt�,N��d�ξP�ߐvޯ5���������lVҟH-����V��0�k�]���I�!`�+W�� ھ[ۋ'O�cI\��e(& ]���b���RAg��&J����Y����f]U���"�ǎwZ���Ks!J�z��n{�.|cJ|��������323S�S�0_߉q��ֺxȐ0�/�Hm��z���A����cnh}���=@R0��u�WX��� <I����K���3�lee�����?���b^YԿ��pG9Ն���P���L(]!+9(\uza*�����}Tj#S:=�D ��g寧-a?o]��[U;��?��K�$��A�	΋f����L��<jX�R��)��=M�i�?U׶}��{���V���CojYv��X�#u���=V&�!)��XU��W�����9Q$�����"�W�`�	p�CcX{e�Ð2��x�j+�3l�b1�{�Y>Ba��ӂo��)ѐ$���3�����~����3|fB��:���ߏ5s~�Sb��КqZxF�VTM��QߴMI]�m��v<o����ce_R�����1J�-�\/ky���Wk�~u�Pdk_Ṡ���SjB�-s#޹�a���s�jES�ͦ)��eR�-_�%����<>���f��vv5�4������Ro�B��M[��0d����ѹ������k��f2ɚeϩlP&�e=څʺ����&8�f��=������G�t��=cIpn�6�V�B�@pF�"sL�N]�8��J��H�Mok�igE�0n��)�b�*A.�B�փc�� sl{��H�!v�ѴΊa0�@��6��jC��U
A�wS��yP�Ͼ(lɪ9�l<9�mT�����N�ܐ�wN!*���ۏ�����/Qb��Y���W�V����B$�K˺��ʙ�V�jX;$V�� � ��^��П�}��ަh��+ѫ���wIx�F�m��=$M��a��b��O�2j�|ml�q���!O�M�|$lMc�p�p�AE��1��������������q	ǘU;X�D�>��٫����f��[��	4G�d7�/�c�$4�"�O��-p����f,�I�v,M�=˾��(�7N�7"8g���R���c8>�wP�塦�L����������{{}MF-�Xc�>>��$i6,J�*�f-/�t��
��!LEl�K���jA�=U���� x�o�O�<��v
)�o���U蜂>�G�I����"�ߟ�����p�q/�N�)'�ۡ�p,d$�E�dr�(f#U�Q;2��\r5b� ��b�0�80�'�h�D=���8�t�Cb��(6��JR�7$���U}��ū���'�f�uT������ʸ�S�"��?M�0��q��;0�a
���=61�QT�T�<��R�^c���ԧe�xU�'�e��x�L*��@����[rc�<ᛜ��&/��F5^ɁZ#W~Ji��jU� �5jS�~@�6�4D49|�����S<��«�*S����F.EuT@E"��C��;ikn���NJ����?�m�>oɱzeRd��/y��`UZ��ȝ��1�Y�w�cF�LP����C��H�:�Ҍ������wS��r�1rW~�>i^T�,�w#\'��ov�c6*�!�λ��ܮX�V�5��R���@����n���������b�V����4��r�`g	L��)�VÚ��ExH&�o�u�d�A����b.�Y�|͈�^:�K��W9v��!Pm�@�<�8{���,Cw�4��?���l�a�,%�lׇB�8�sz��[��Ƶ������hﳇ`9�zL��J|"G�h��>�]�1��QZ$д�gt+ɗ�)Yx��`���H><�Z\�u���Vv�]�ވ��B<����T�>�?��\��W���ӬT����2se��S�ʍ�uE"5��*HF�L��!��6>o��~���M������(��f�4C�/,�Ü_0�[�c����u�X��0LS)�>=X���p�y�mx�������:v!���a�S\����hzrS�5L���A��Q�Nm�U�4�y�F#3�sEi}��]�l�,�j߫�V~�$��W7~V�e�X��}�:��W.�����y��R��q'���N�C?L��/�kυ�+3~�dN�ŀ�B�zF0|�4�d��~���A9�i��䞬���#������wfQ������5����?Tu��-����#����3ﲥD�7���@?!:f0x �).� ���L�/��������S9����>Rw���b��n��i��N��5ɾ�W��S�oy��PT����#���U��r"��]��釭�O��ڊ�R��"�D.���3g�2�����pJ�N��%W���϶y��F����Yd4o>_w��-��邈%f���r�QY�)�-ʿ!Ϊ�^��A����|��a�C2�K#��Ĩq�Pd���6���J���/��Ҡoxy��[)P!��:m��	�s=RShyb�� gd���C;�?O�h���Lce��"�nc�jCM��zz���-vy�]��-2���dk���a�ZJƎ������B٢r�݋q���=t�Of�� �)RC�Hf�pV%�F?H�벗�f���?/NV�9N�Ы��~,�<���4�z�3o���D�����9�P6�I����|�k;�>�������VE��i!���m�z\��M�j�un+�����An�ũ���׺�e�`�S�*�I��\��v�z����x�|����04�am"6�=
�,IY���ex��N�������ځx�4�)'�3 !۝H�b�(�`��Yc�<�%�P^��7xӬ\8WrK��ga`\���P�Te�2��#�#�)��%��ڃ䞎�S1:�@��	���)"^d�N��j�^����N8;  c�q���&�U�8��;&�km�S�L5�sB˭�'L�|,F|a�R|U�� N�a��	CѷWȁoT�6���XXn/?u�ݖ˚���6��8�����r�lf��̾~Cf��=j�'~r�p#EC���a�t�_��wy�9�t�c����MJ[	nY��`�VJ(�������s�=�v�N5I�X���1�ю���ý�̟��15K�-Ɇ\yx�i�o����ٙ�E]	r��8�Fݍ�:��V�_O�3xJS�'i=Q��D��P�Tk���1�0��xM,�������,�A�r�=T1�H�F�-�?FC��Q���i5�2�P����O�3�� ��@9��po�N'k�!����ǒRt�c�)�]�镼�_���9k�֝yCv�VO!��[���`~��nf7����3+W;o���7��O���yW��of�b���E��8X����Y�/Hoy���ۘ�x'炐E-
�,�-���ꏓ$��,r�h���}�vZ�֤f��"��' �,xeQ�pz�e�ɿ.��g+�����R�ȴJ'1(����mn��8������E)^��@Hj��2���)9O��g���ʢ��Ӡ,�������yK���1'`�Kظ[��y���1Xb��O:&J�tlK6��B[�h�*�4�.H�3��f.�G�Ħ�*��%�� q,�v�,������->��NSp�O�����}���b�t�dߕ:@�L��f<�C�Om�r@E�]�\�`����a��t�+�j���;F�Gzz�XS�l�Ze11�J1�Q���;;��Yu��$񒦨`"�9�5��x�+��A>`o���/ӅhBH���G�O������qT5�2
,���l7���~$�e:��z'���ʍ�R"`�?P�p�	ev�"�GA��|#�cs'rd���ԭ1Tե���86�����1f��xX]OS���_V�f�:{r�}Ӯ�����p����"�`Ոw�fn��"�������/���:�����^ȭn�|��+<�V���ә�o����b6x����)xy�;ˑO\V��9��cQ�yZ'0	+�~�����m;�7�+#-���!��0�>I8h�����JeT�<"�V���~��:���h�2Ƅ�&GLh�����/����2��]	,v�������Y��@�QbH1W�H@��%;<]���<�{d~�"��.�w���Jf�s�r�7A@Kto0@�`���w'c�qK�ͣBL�Ŭ�A4�B"-��P��!�~�!Axp$�[9[Y;��V��h��X�>2!�v�y��N&*��_���b:��oZ��A�3���k&/�������N@Q���]8�k��,��j�#_M����װ"�w���1��VM����U�ӵ~�4��K5[6�
	�|��~�Iq�X��TP���v_�S���}�6ۙ���Q������q��@Sn[m��7B��2)���Y�fq� w%y]sR�q.�B���"���W���·��e��	��$ п!�E'���2Y:����<׎���4������oa�}�b�Ο���QBՉ�G����Fg~�Q�ȥE��d)4�G��<��wR&��w!4�
�dF���(Y��W6Ů�(���]�D6O;bs�(���eM�h05�[\?��h�F	�-#(r�yB��1IƑ����t�?G�ހ�~�:����.��{;���� 7��L�o����y\�( q�4��o�WHS�O��h�AW��Dɕ���� �l�ݒ� sF:!��u�0�W�d��>b��*c��F!=�@���V�n�F�4a�T$����Le}�v6P[�ʼ�"k�ո��oE�O`б���Mo:&ˍ5�:�"?5݅���5`��^cv����"�y@6��t]�Fh�D���MW���*�p�v��V�!��^��rf���1��d��ns�C?�&AT�&�d���ҕ�k8�vXi��R;@0�%a^��o��-��K�sH������u!���,6�u��iTO�)��~��]��M���n�+�+r+#c1�W0��J$�/?�A�n��y����ց�9Uﯫ-���>��\ -�w��v��%*�ď�`@��������k�O���7�&�=j�V�JGmR��H�˩ly�z��ʳ��l�����\	�v~�G�id5��0����
��g�2�(^~�L&��vW[ke����s9k؍o�{�A����;����".˴[	�An�I)SO:)���N��+��neyy�d�qZī!�; +ϜnΒ{Sؗ ��R+�	�򎽜�I�J���d��n�K"C xiMΠV�-�q��d��@���0 �d�sǏuB��C�������?tE�K��`NJI��JnĶ��k*np��HM�T�y�9{�L���Yp��e ��1.K������S�d6����P	�ۼ�Kc��ѐ�LV�ʍ"k�]��`d������وy5Y^QOR�d�����H(O+�6(�	�#0{F`�i�6�SYJSv4����lB/g�˿�,��K Z�o��Z��2S$F߼r7���.���TQI��3���ϱ0�Rk��,�cB����;���ځ/�^�ŧǿ��:�i_�rg�[U���#��=(HR��4dS1OmlZA�	�V��ի��b�\��p�^�a�V��p͝,�aԏ(BD,j�	���������m69�-ӌG�OՄ=�A��y��,#*���H�+��Zkqa�4�n(�!��	����q�ǻ�{�O���2;���z!�U�G��kn�?Y�T�����6+���k� FV���@��~���xW�����=���f� �)�aX�˥jv���T��r8�u>��48��:H4��	���t��ŕ���{�la�<�{�HO�8�ǉ@��Ю��R��8	rEO�)�?���-J���/,��V����f.h�f�7ߝ�{#r��y!��,�>�B�`䙶���Z�l��x,C�/��}oi�_�>@=mt�!h�n0͊{��IoT��n��²�*M:�jW_��2r�r�K��1��ev�ߕ�C�w6��MS	���<�۫��(��4򼟫�D�T�b&Y�����$Mg�$մZ驆��X����ێF� d%,;h�*->�Ȭ��%V>�S�A�X��>_V�Q7��R6�o>�� �(�oi���h'��ur�ق�y^Au�Y3W�2��Q����i��0��A� �dZdf LNk�l+�%��{�5Mo����-D�8�J�b�q����K����o�}�}EF	#tG�3XH��C	��������ZdC37��/���m��y@T_G[w�����cծ�\9�]���p=yԨ0����k�n�>b=��䣊I8X�%�߰*N(��O�
��V�7��F�wy
˹��c�>?xOl���6v�|zl5e/Z@{���:�W|��B�Q�n�����r�,���G
{QA��FP�L��*�i�,e�O�X�`$��df:��7�jw��|ߐy>Q#Β����$[{d0�m�B�nT�����lG�{�E����C���N�:	{�#+Q��6/C	�I�R�b���ͧ.���"��ԭ�a��L2(�.��bmFT�i'}��Gh�U�"r�ǙQGe;X�怲̔s��x|�xHf���l`!��<���#Js����K�����^�~�E��X��[⦞кN�(�,v��%L/<J�@[�b�,wT�)��H�����66��x���Ȍ42��N�d,,5�_+%�i�5�X�%����)c���9/�_k択��#il��k�.FJ[`��
Vi���ަ�GM�������eaz�*��T���z�%��y�.��<���Ԩ5�E؍IX��SϾ�Ĺ��x?g+ޒ�I��:˟V�Wp8	�V>>���\��ddJ�����s�E@�v�jt���=�M�;O5�d�����c�4ҫ������q����76�Y�fl�9�_��4j�vb]6���� �A�����I�qOK�&��S��l^��)t��}�C�?wfI����m~���r/ng�ꨟ ��o_tt�'�&l�����4���(�Tr���2@�U\��ano��κ��,q�7Ӗ=�g��}G�0,Pa��1>�Y�W_���}��L�3��ć��
�HH���4;�L_�֝E~1֭����)k��1�Y�W�?4aK��k�r�$�?��^�sGg�(�8^�s�2��2q��|�
��E7Y:���b~Aew��|[R��mD��6N{���X�*x��y;�C����@^Pv�#.e�_����"N�R3v�c���?���ѷ�z�d��0N`C���M�K��t:t3z!����0�½����`%H	��M�ሪYRL*G�ezT7I܍��?�/c���L"����{���P5փ�C8������?EQS�L���`�h�0�0exD��] 缘�kf6e�-���P��� ;m��o"'��l�� �+	K\�cD��{��!G��atf�K�a�:�5GK���;����8��s�9�d��+��9CN�s�����ZHD.�IN��ɺ�h�I�JJ[�hG�<:P5ݏ�Ӓ�T���N_D����s�;�h\��6��i��ư�=m��]�r�t};�v��p���]w�q�,sQ�	ꃛ�̀�o&QQ�J=��(�j1�����wA����7�ի=ep�8L����5�&}�~����M���ԓ���6Dlt��3�h{���倿@g�
P' �������8{��a��gDQ����%�z@����^]~��������b�MH�)�j���*���+$��[&�;o�����,��grZ$��}�Oq��(.V��:��j���1V�N��.����L<��k�DDƺ4F�8j>yI����p�c��D2���bFf��[�3��h�]�[���G��ē��2b7� bm�����ٴ� j	dbৼ�~N]2t��~���d ���t�X���W�;���/lz�s����xV��p�)2�TQꎛ�S� ��鑾'ٕ����E����nW�h�a\6[+��ד��1�����w0����'�2����-��Y�gl���tE���x�d�wv�?�Ӏ�h�����2$��,>�Y�Q�ɨ'&�$���������m&���/���*��!њ�Ě������LA�4u�WX���臨ĩ��Խ�=���9�X�DET�ն�H��rBb?,kr5W5ë�9��M Z�
c����9G�],~���S�=ؼ\���/<�C�x��x�\LDŠ-���m��ac�����O��A!�F�E=�Ȕ+]z���A+o逍 �ӡ#o�<wZ�T)��'K�yE�7Ν3������l�r
�,R�@�]��#�~� 0r�5$�V�v[��\����ۮM�U�/��Mg4�Vކ�.n�t�����*�j�n*zFd7d���X�o��w)y�$<�yM1^.�(�T�x�ľ5wx�f�,xKR'N��W�74H\�}�'�4���2�'],<M��'���|�&�����v�?7���RN=�d}�P;B�����C��O%�4twg��w&��J�b���zR2��pٵi��i�t�4�,�ïD(�	��1�����ϲ%���m8�9��f�o����4 T�3TVI|p�r.���e>`�EbK���U�i]�a�"M�iU}Y}#��]����ˊLa\��uN髱(i9kdCw˺Mv��s�"	��Z:P ���+����b:3ax����Rp���J
 ��|9����(�dÌ��1_�QL�[_�@޽ ,�;��YE_x,��s��Y��GL���RWC
�fa".(�4giK���Lx��f��Sb:�@�� �HQ�x"<Z�4���%ӭ�'7� �sW����缜���,EP�^Vx��D��6[46�H�V,�@��=۰k2��"�~�i��Y]wx]ti֩j�́C><ڵ����gj[�
(A��P��#E��W����-�	b4�4p������o)J���&m����UpN�N���o<�
w&���ȏ��纉'B�,�9x&�'�s�:ǚ����=���xtdIQ�o�В߃�/\��2}?�C}qq���n�	5	�y}�|�JRS�LB�z��ȫ��7���l����2Rq����I�W�'��¿yU�O��k�hf� �+�9��d wu;�.;޽`6\������o�ϗ�Gn�0��{��K��h#>U�R!%���Qr/
��wb�s4Yd"R�_	d-�0��I�Ǫt�V�Ǵ|�ֵ��~��jz�2�-�8W�� cU��5��u�Q=l�]�W2�)���XEXT���,"ǼI�*M"�����jm�2�LN�imU#�IE<�1���+U�,�~��sJm	�aR��!V6���4��G^9���6���i�Cޓ6o�ƃ�KV�(,�(,���e�Ǥ/>h/m��,�Ϯ<͉qs N���ŷ^Vt�,$wζ�s��x��.��a���H���4����pH�h*v�r��y�Ո�j3��]�-������(�L�u�����:M����.�?_Q�����fuT�A�.&U����_I�2�Y{6g�������~ x�C@b��<��D��K���od�,��^!oխ.�����@Hc`���c�NRN<e	>����4��pvrW�-����[��Rń/2�]�RR�ƣZgq�:�[����\��vO��`R����vH�[M}��6�B{P��z�I�O�g!`;�ƷkfV�S#Ww��od;�݀���uɎ!�<��6#�2A^�(���0^q�ػ��C5�:c�x1a���8$)-�zǫȼ�ٌ�h���Y2�Y(c�B?�#L�pF.:��zS$XS���
�������E��ۯZ?t��r�����C?�Y9��R�O߲D��`�c��
�]:�f���~����	���ʿZfaSf���%)�=�|E�P�-���TqWc�z�n�g�%Ϟ�Z!h#���vN}쥕t;��5�`3Y+Q9."^���2Et:���]FY�?�1�}|�v��Xl�B���kn����u�m@-�#����B Ũ�V�se6lQ���	6���@�jn)�syU+_��i8���WUw2�j�/����Ś��"�������S�ύ���򅭩Ɍe�Ѝ����@��5I����~�dF�+�W�h'�;l��^<] !F�v��PA�{k�Y�1���)5e����I��(q����ʄ��Q3�I�3ԁ�#�*�%���O�~r�T��w#C9�j�f�.�f�C:��o��
�������#���n��^��F�l�ciwCE����f[D�[����}���6r��e�8R����!$��9ѝ���.�|��ς� U@���^��T4
���m���ʆ�GFZ瓬��u�}��"(R'T�����nNDF#�a�ӷ]�kZ����o�ٕ3�H��6�')i}jm�?� �|
y�*� ���#������Ag��Jy�M����&�r��a[��a���[3��j������^��̾*�i?m�$nD��^㘓�D"<[t�	�{�@�=}�?�w��K���`��Ϩ:�s�E@[�jkt���}��;:��_+ I!�n� �Dm7�dM8�(V��c+dήF��f�����UU�ѧ�HDHkӜ��-����!���r�>_�FZ��Rp�J�f��1n���g�$��.�5z�#7/o��P�]l��E�+�U[��e
�Ц�XTV'�u���K�2:V�K������<�+s��>�ޕ	V�R�2��X�8�F2
.�d�C<�cVҧ������*خ�Ob7Y�M���j��l<J��n�aDK!�5��u�{�m��)Ձ{pu�X�;�L��� ��3،_q��Zɀ^���fq�m��$y��/"d�IQ�����M���ir��(Ϥ�d f�|Ty�������ݓL.�a`έB�)0hw���0�ٖ?h�,��R�Lt�7��7��ff�t�#���CEc"*
<��L���@��4���9)9�)?���3���Ⅾ?(��ư/��QRSj��IA�Dg�Fc�+���V8�������z�O}���a4Ul4@�m �x�>�	f�4�M���J�-��r�򟲭�d"P_��?�g)��7��~Q���ë�F%�.�gYή��g��=�U�e�xDH�D����3:��D����':���PP2D[+4�J;[}�S�&tMv�[�)+u����-�Y�ȧ��q^�Q��k�����a��6��O|��Y�gRzyTL�YN����1�O,�P2�m�>B�{>�UU>�&
�M8v�֏��t�_��[0�v5��u�8�]����]��?�	�����,���������!��A|�,��� ���TgӇ��" �����kS,Uyʞ0w��#������'�4���	��Ց��}z��0L�ɑ�DD�*_=#�s=�!�8��#1�)�	=7)������\���,|AN;O���܆wN���D��09�@3s��9}OHcI�c�|�zzU&|oB}!�4��6_#�@��4��P|`�t�$�7�ab�(!��v�
]b��{t��7�u�]EJy�_Ɏ��1��Ab���ț��:G�ư�y/Mj<�6����q
�q���Vc��$|��O�%t�g��"�^���/� �P���L�� 3T�҃���~��� :׻f��r9l1l��b���Ţ���ܧ��l]R,�5�(c�m��&��s�^bf�����j}q���Nbj7�Y���Z��\69�/��jQ��A)��j���WQ���K�σM���� .
���:&�U���C���Аs�2j{<H&j���y���w+�<���n���_�>& �Cb�f����aj�G��X5j,=ݒ�o��iOJ�.�Cj�d�|0�����nR%�%~<<v(��hMAf:.��lL��FX�F���jJsHYJ�h����L,Y70�x��
��H�X#/T��x!q'��ſ�<l��6,s�BJ�E"P�(�� ��i�+j<���������, ���x)�v�8rC�5Bpi;c^�>�#�t蜊����a&�lx�������o���iu�Bt'!����O�)��|_U\1 �㹂&J�AR���`fI�zx�<ݨ�S���Na-��5M�8F?�$T����t�EV�r�?_i[�^�ׂ-H��4&���	X�t�.M�>]�  ��iБ�A�\�y�^3��U��G)�>�����w����C�XD�ɑ|K��(���������wO�I�b��N��/�d�瀙�^��í8��ڒG��x��3C~5�@�=��ؾ.1}sb��s�iA��k��n�DUMJ�1�ɥ�Q��rbHG��n�B0YO�B��Xt�+���6`U{k�f����P�%s�Q]Ģ0X����O�K~���H��*}D\?���W��)��@��B����*�RB4#��"�'	Oz�ԽȾ[�����(UT�V��ʃ�ec�G��U��J �s�,�@�|�K�YTL���)�d��]�ۼX&F�v}���Ie.
a���2S���SY��:eT9��G/-V��*>_� JM�5�e}�'�~������B'�����V��C�4����qco0��,���UDX�d~s�m�����LΩqP��2���hm��������R�ɨh>�@�2�V�����p�(V�~�H���<e;sA���Wc'W�I���R"
~�`���>�
���Z�;����L��cu��`5ͨ�d��'�x�n¼��,�ƹr�!y�'Y+��чl�U���ј��L:M���0Nt�#�dJQ��#�T
K� *�S�A m�DU�r���.��в��@/_������£����B#���)xbk�a;�j��;m��Y����7��%����F	�e��BN�0�DU7wqex~��=�C�27�KO�>�t<0OM��=�?B��<�'���g��> �Y����N
w*;�B�d�#$���Q�
�B����F(�*��B]7��L9����U���`������:KT��Dj�	�Gq��|�.�:�d��� ��U��	��i����9[�,iH��u��<ѓ�c������!�i*��xđK1��|$H�A����8ue�5��	�.J֓k������F��