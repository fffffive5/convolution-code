��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<���I�����&��p_.��㥶��<yX�6���@+R����;�sg�v�-���sk��%�K���P�ڽb}*�pQZ����O5g�/���*.]@����o��4�����Sb3�-#)/=p�`�_�c�:�dh�_:+�#�׻�p��??�F���(��Ac����r|�Y����/G��C)*�d`�x�k������
�u}Fa�yp;�����L1��o����y��r�%m-3��<{��d9���a��$��"g��'�6�@H����cm�8�3��[�$����p�g���qqDj@e���X��z-��hK_�c}ZM�%N9}՗0>�!�J`/�#�YDe�
1��k�Xz����|hNul.vḏ�A0��d����?4��@��{�R������(�5U�g���2#i�S*��.�G@��݉Äi/g���]ѡ�����(��ߨv��l,��䑙��%��
�>P����H[!�_aw���E�d����z���w��d$fXYz./�\�T�LR�����u�$��~=*�>t� r�]�0�ə�}:kӤ�͡81u�*z���a@!�����>������E�����sf�}�:�ZD���l�]*!̊�av~���j��t�[݌u߁��-�F`E���MR��e��]�;i˝7g���l��@���C�z`aZ	a�]/�Q�*7b�Q�/�� ��1�����\e��&{�ѳ �\�5���U�������v���wgi�VK��l'�Z��`���6�x��:�D�/�m� ����X� ��F����ܾ�{~&�>.*��]uHZq*���g>�$��K�NU��l�A����������ŋ�k0�h��/������d �g��`�Fg\ax){t+gT��)Qc�nD��ͣ�R��K�8�k�E��]�;�������E>����$u�m��Yw{XP�VB�9��1%���
f��.m��A��k)���k�܂�F���_�ph���j�Ś=�`Cc��P�1�J<��6&��.��K�����&�$����� ��/�mmtikwc^;�bI�PJmɁ{��/�j]5�w�	H��g�%�̒�����b-]��p�j��o�.{����t��/����g��rU"��^-�]��&	H=6�OƟ���k�Ge���E���������+o.��g���oF����՛��5?�T����d+?�R�=��A��wJ9��+�S�sjQ_0r���L8!Kz��y���&$R��j��B����A��3�wA��z�8�ztɺ��e�ȓ���$�S�(B���T����ԧv �ab��M\����QĻSQ`�O <����<���'z��-��Ę���R<0�k¼�IH��El%Lљҟ�*�6�"�NPuYY��f���T V��oB�Y�(s2��, �"��!0�5���Vu�᮳�����v0S�˒/�I��9�?:+�A7�skL^O?��m�S�n� x���R�'���Jso�q�py9+ܣ&;^}]ȳk��%��$��>�А(���0��f���tS�pf��B
�	j)�]��$�J�P�ɦ|��d� }h3�2��}�!.c�v*���s�_��D)��ۓ�7V^�Z�U�g-����7N�u�¡�H�.��M��ue�lE@��V�\��Z=��j�OhV2gju��s�x���W%}��`�a�����:4[x�5���r�)%z��]�]!p��A��Ȼ����
cg��ΐ��`��f`�7U��%�YeŊ0$a�paX��W�ȮB� -���J*��éKC�$kQ��0⠙�a�U���&�~�j�l�r�ؾ�~y�#��U\b�&9�_f́����Vp��C��R@K�a5 H�t�Z�`V;@��R�t�[�|��A�����7��9���xx�%�����0Li�"�.����{�����"���&m&��[_�61�����9b�u뻺��H�