��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<����o��t�w�H���vG���lk\�~�N'����P@�����=(W��u�:W	�	�ț�:��ɕ�h� �8w+���f������"\M�,�Fi��������{�fAٕ8޳�����m��o[|]Ԓ��,�p����~������ :4�y��rK)#*�C������6eʈ�r�t���	A,��Pچ=G̤B�o}�F�H{+�.��qɲ����5O{�4���"�J�y��LѽV�q�~����e�t����8Ƒ�L����u6NF.��>3�b�M���XkȽ�.�Hd>o�Bd�Y�8�p�$�����<����yS�2C����a%��m�zJI�޶a|,�B�����N�E��p�\����F||��z+BY���90UA.�辍pl
��+xz�# ���%Rvsq	+�\5^3,q�V�fބ�\=�Q�/0��9�z��̉s���@�
�xd�_�J�ƃᄠ{� a��O@Z�m, ��>Bi���,�y�Й��<�� k���������F��2FfC�Q=��Ǘs��P�Q�B�1��8�����D�g�בAa�M�tʋ+�K��,?؂1�%���ŤF̥t%�|[�BM����&�� ;z����O���]�Q!�ofv(���؍{a,im����/֨9��;؝�>���I]����*������ �w�msp�@���B�&��s<�HQ�ăK!Ŕ�Ok��i3kGq<�-��7ۅ��Ax�aaU��r��r.K0�n��/n���(<��Pأ�㮝Tw���M58��G3���>�K�B�mIq����1�|�E��������	��*�i��x��,!�~��)Ӻ�aU���P�d�X��u��M� `n��W%�Y�g�t=mKR_�Z���ݨZ�����VE�&ߺ���(M��e��S� ��?�܏,��jQ��0��nrEJL��G���/S�L��i\���옟.P���K�q����;X��j��_�����0�Q�����Y'y�b���i�ǚ�Rg .�����~j��
� |b����_Ǹ�,�m��g}?���m�.��"D����#��q_Wy�3������H��~F��A;�u���{��nK������=<k%}��GU:���[ֻp4�X��,�O�CK�,�D'�7*��R$E��0c�$b@E����Er��Z���S"hmLZ:I��=�Uɣ����+MDK����n5�;!��Ϛ�eW�ڡ�T�2&K�Q#��ߢz	�ƒ�.���P9�߲grg@L���)���b�����p�^|Y�{J��(o��T��h$���*��#�S�ym�K�}�!�����[)��q�1U��@��
����G��bs��������-�R�"�%t|�ՙ�UI�R/ע6QD~��F�2y��s�w��&BО�w���	vÛ�2m�:�5=jJ6@�n�)%�/�%\��amݗ���J9F,����-���8ʓV,?��C�&�l�wl\HkKPy��O�a��`
�ՙ�h��F@�,D���m��n[�Th~����s�w&3�������Ό��p�x��cK��\����GT>�h��6Hz?�Xk.w�St���r]�9�̮�d�{�e�`��%�ͤ�$�$z���|-ƴ�@|"D|�"�D�&dc�T�� ��������$ ��;~E��٬K���6@�:%碥�N]�?�N8�Q$����|ʐ�.�f��Q;�^�*���/]�C��U6$�t��q��ٌ���J��̯�~Xҝ̆���^-YÑ��Mx��U�O Yk-紶D����-N�ZmB_Lh�HB�6�'6�n�hk��JI��J.%5Q��(�:�ث���������˂lﯙHa�X~HΟOm�_�U�p��H�B�W�$h�~Rw|��!��~;<���^���%b'}���^��k� mDU������9_�S� �����B/k�7�li�51;�YpU	�}"�R���(&J��9�h��A8Y�H:�B�E����9���$ܤ��C�Ha[�`�}� \n���R��n/ܟ�{I��#�!o��PZ�^��y�����	��Q=���/�/�����	û���5�h���`�̨ y	,h7G�+#R��ne`ې2ځK�e�_ՐE�ca����Qq�sR�朧d�$G�Zh����,�Pz�:e׀_�!��'z�'��|&Qڌ��i ,���|��`���3
�n���L�򺾲�?�rhf��\�f�Z�:���k1��� =���D�7W�oy�#>��,�u�~�~��b�K�_�u������<�B+*M�iGv=�1t�^��(h�1D��֌�^}r�&�!�Ѥfi��q���^M-/�^��+�5,�rE6�ﶴk���*X?:���R|�ӕ��͵{�Y]�26���<�p�e b��������>��ۢDs���}�#�`|q5?�~�2���Q�C��O������� E.�0��G��/��D���O]�����Rob&�8څo����pF���bIu�����n�'�VM�����dɉ����)7@~�a�T����V$qO�1�ϐ���3��uY��V�@b$�&�ʎ�&xBSՇ������d�Ч���.k67��R�Z0���:9����zA0��Fkd E	����ߵrY�B�q~�*D����yFx���1?ȏ�؆V��O,�Q4��U4/(��� �U�^h����six����|V�Lo+�'�{܏��cj� �HNdh��-}B�20Q��U�0}�R(j�1>��ب�-���z�f�8A��{��<��Y��_�8�<h�g%����5��ڏP���L���8en#�#�$V�ͻ�9BMu���$�r�����zH�T�>�c7?��On��N���=H�}-Տ`6�7��?z�P���G7��>5�� k��� ��B�32���f,�tBu����ߢ'�&�÷P��?����Ht�Y�b� ��}�%�qG��$+K�g7����x��̳���m��m��=?�6V"J$��Pgad�*5 -߬�J���q"Pm�Q�`|���1��¾����r�����J綧��Z�:2�=u/ǥK,���5{	����#�C�_e:� A���V���;��r6���X�`�h�dUN���