��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<���t��ej$�	��PiC8�;��;������RR��Fl|�8!��<��_σ<�;)'yW�78�=��@ �(��W�Y�A���t,#^�y����"q�$}v5X����^����U,�%'���ZK�`�X��0���[Ԩ��L�Ɏ1�Z�Z�`�P«���J�]�ac���on։ft�2ZR_��'>'� %*<f����J�Od�<��KD�@���"���G���3������E(�Ρ%�>�o�=r�4�*���X�w�#���/�=KX�{����z5"���U�w���:�=1���/G��x�P!�$���kِimJ<��e0�VNK=�} �v��ݺ� 	��.�,�E9*A�kB�cE��o2h{'�@�7����S��@������S]n���ݟ�Xt�IxWȠ�1P�+P���X��<�$�c�U�B���*���/��b����af��������� o�{��s^����"@lx;Z������{�1p8{�%��4:��@�;���g�u���;������=�"�Y�%�6B�:�F���*�C��>��%c�Z2����zo�	M�I����k�(��^���A�~s��Hª��M3���T
�����ᄉg��MBHO^�i�"g=�t�ׂ�H�O>j�ɲ�n�z�-W���=K����١�38�I8R�i@JlNn �ӽU�v�-Tyml�P�S�̛��Mb�r���o~`I]���Ǌ��6jN��[5����l��D ��P��
�_X�ʽ�M!n��cK��Ƶ�NJ�e�{�����
�LS�L��TWQA ��Q��;��F�{���I���!� ��n�����i��;���6]����T����������>�A��!���e��nB��Q�r�{��~( ���s���J�i�{�i�aT�n�)�2 P����@����K\��j��~�EYd:Q .'I��Ҋt��b�\d�k��������eqpS4�Jq���c^�/�n4Oe](����v�I�_C�3`)��R� QB'�v�Q{Cl�d6��X����,�IG;��>k��c?��e-:��i���[~�mIV�n�u�y]���?0Wt���uq�/7�ƥ��MëB��zφ��?��4�'�|�v���㤮{-�=�Y������"��#K�p���
���pc��T�(v������?�usD�O)'���]������x+e��@���@�ꕜߗ�s$�8mXC�"�C�e�w�J�:�{�ڳ�,g՚Ӭ������_�z�D&-w�L��D�9<0oq��Xͽ�����9��&�W���5�Z��0�;Ϥ��@J��~�ҽ5�ql��r�Nv�� $���
��=�ާJ�7�b�O���d�'ñ�%���㈊	X$A:�M��C�~9���'��������!ȏ(�޷s� 1)��lSBx<��eH�̀��i�q�WjuK�S7�~�cJcJE0������^�A�U� -?�5�j�����>5�34�M�k?7#_<і枑��,�t�����S{�uy�ga^B-��o�^�0.���$�����t� ǋ��}�gWC��LI�Z��Q�a�e�,/���m�_��@�~*<��zȸM?�	7���ҟ�86��*-؊�h<����ޝ���oP�u����q��U5��&�Pne�ӓ���r
TИ�J5��D�k	�)i��� X	�n� �~3�9��eum��҈��c"�G�ܚ�nI����Û�y��nѹ� r`�?�t\k�/a�B�Nr�]����t�vp���_�;}G朂q]���R�sg�H�B����&�pg:]�s!�x�}��F�6��-���8���2$�EA�p�i؆�|����]u����?����53r��{Q����c��ˑ����x�J��*�(=�H�Ƕa%>�aId7�TX��ٝ�4���ٝ7���kN}Gu�8�����1�4�|"��<���;&���ӛ�3�؊7'�{v�F!Eyi�:]7���N���+�Mo"#C�-6��¼���\KA*��L�t�x'��m�L�3�4g���V�v���ln6]*���Q�e�nkv�^�dbK���E�ZG;��:*z���$��C�ƭ�x�>~��ÖS�n��$�s`�����o8���
k���S�_�ڢ�|R69����`{m��y�y��Ǹ�
�?����i�2�Wm0�:a�Q��CCnYى,`B��社�LL�}ܰ�$GE��:~l��1��/�Y����јys�+�f�p���l���\�oʏG��7�:I��{ߌ#����ٯZ�P��6��T"���/p���L`��r�EV㩼p�F$]s��F{z���;���#���A�
wT���8�8)��q�.�%�Uv$���7��߾�RN
E�6�f�W�3
4�z��)$b�]*�$�51g����]�*N����̣7��/R��5(���;�i3ݸ��A��2Ka�f!M�����2��&n��j�9�W�;ӫ0LX��p*�fb*������f���Q�ƃj1�h'n�ϯ�i�C��=�k2�|�&�����^p߿����,�y"܉���4�/��O�JB�J���
��� l�Li���i���!��T���X��1v��@T��1��9}<��^G{�g"�YV�E����v��-7�n��,/S��w�|2�S~T�y4��'Xl�u"���D*躹�d)yd�ڨ ��n�:.�
�G�����T,��S����	j2��o���`�+���a%�\;8ৌ�v�ʎp/k|��Ӂ#L���Q��]ӈ������lWC	�ٜ�j�W2��loM9�6��(�:l��c��U�x�'��p hG�J�h�h�T���k�[՛�����S!�;�.*��C���utyc�[�E��x�#�q@��:��/�����q؆��a�Rm�mEN�Ѯ�a���{���K\v=����	 �DHET�sR�E��P�(�-��f%ߴ�ꎈ�]�M�� ��f��B��#y�� �D��yE��T8F_�ݴ������#��u��@_��#D�S�#�<nZ3��-��1�� $iIJ.,C1ٱ�q&N`S	C#P��_*�S�-e}�V8n�8y��������zS��+��Nxz�c� \I��Y���ݫ������h}�'�R%���A����2w��罻:�l���<��9ɵ�0�z@��"}?DQT�������ɑ�k5M�9:"�Q��Iq�9��Ԗx�!����W@��gas�Bާ_�;�h;'aq�ճD�fc�����J��ǑG�^��m)3������9YI'�*ȥ�� 	sO��Բ@W���
��/B`B���:�w��N�e���U5oS�>1��I?d�i��n+� S�����}�Gۄ�mr豏*E~z8�_%��$�
㹅�,���V�����I�4Q�
�YUK}��k�H��oA��}(�����C�aoP�ǔgr��f&�v���kT&���7DwH�\��{PR������U-�r�h��[�o�{ �����ʫ m�Qp6�XA�@�h������"�F:̼a;;���
�pc1p)m��y,J�
~���{��.�����#�C�L�N)9G��k�D�]�p�ػ��v��1K���C<b?�^y�s�(2���$�4{�90n�U'\��m�8.�se��\��{K�]uZH�}X�5Y��*F�q�z��+��s��;B e��I�B��6�.��E��'�U�����X�ߵKwZz�e�y+ W6���?����uF&���e�ha6/�j:�5-A�v�Ǔ�@J�[��'=�m��7<�Q�u#a��e��P�aE����Q�7�UⱠ�3TBa(#	� �������cZy�&,!c�b�_P|ޓ�p%���,:U�(ұ]\�.	�yD�rτ4�Dȣ�I2!���d�ތFt���tk�+0"��J`�F�c���K�����
�:��e��)
�pRN9˺^��|��	�b9T�gZ�{�OP�����!��2�Դ�����S$�)q8~�r[j��'`�	}�HQ���D�[g���vP���R�O!�p��e����紵ә�v�����o�o=tT���?��7D�0	����MQ	��V��q��4]��?��A��5|p�Ǿ2�x���'­E!���j�������;G@�
X��݃��(�n.v�W\-[���}�+��]�A~���۩3��Y�]� *@	 t�6v�˩n|,��p@6ܥ�7�U����p�~BW�aj[����BI�)�ָ��h�P������h���X��x�G9� !�*N`
Lo��s5a���
�.��"X�V�h��;��:
aPR	�L�\e��S���x�C)��>b���i�������Zp)i����Ӗ��U7̇�]�]]o�Η�SţM� bH���N�Z�{��v�t�e�M�8;T��g� ��fq[v����LZB����#QV����
$��Q�$�|�s�����V_鉴n�aUW�ڀ`rl����].��Ҽ�޸l��6;���KH���q.�N�F�Ü�yÖWn��X�<��B��,�97d��$#tĜ�(K;�VgQ��!^��i��#M�:0�L�>�O�u2��n�n�2I�4�v����2?m����lN��g��B���<öplDF=�s���� �Ҿ���/�=����"њGӀptŽncG�V�e����1n� ������/&ȃ���p3Ĵ�����+����ZAxB�L��,�+-Rs�$�(ŧ�����1�n���=V���쟩ϐ��a��4�,���.;�����U��z�f9"�̂�1��v�m�M"�F�sHzZ*�����?v����y�����s:��+qwF��f������!�Xs[�������b�D��T#��PO�!c�9�;�$k��Ku�'����-�3C�N�z��s��A7="IYG����vՁ���4�9~&JU����z�Q���`đ5In=u�#UZ���Aޛ�[�<�[��y~�4�<��Vp[*��{�޿bhj�~�wvq���\j
{ 럞�g3"��0&�`���5�����0���?��j�0B`5��9�AR0+������mC�gS2���!_�\%�P�z����Zʹ����Vub?`�iM����FF�����B�fuyj�\���o���k?����=���f�W[CA8%��V��*��Z7S��<�oi��#��{i�>l���;�-�Єp�����3�%av��
�����ٰ�3P���FG��#(�<���@��̌Z�_ˢt�Rs��t�FW#v��YQF�!���O����8ͪ��3��e��B�XUr�#^m����1&Bk�7 ���m(�����3  �Ă���Z�=e�\�I�	�/d01�����ZNVl��T݆䩥����٘ݷ4�	�@V�#�p"P��N�i�.I������*m+��^#�@���L8��	Zv �ݰ��wA���E��0+v}~�t��$[W,q۱�lJ\�=Fƚ�?����h|�7�vU�~>!��	�7\T�`�w���1��vM+l�oȶ��d���^�,#�n���p�R1���:�;��鶍l6V���}�X��Z���Q�^7`��hp2X�
�}7p�:Ag6�[��0Q��.�EdP�fָ+#����
��u����|�= 8P����5MJi@��`$*@)��j�h���!�&�	�>*XR�|��~!=S��n����g�S�i �X������D�Qǁ[�i�fN�H�px������]&XJ�C�.����A�i'ɭڷO}�0�Y�w���X� 1>(|#X�8O��ė�Y W��
e�. ��I@�qD�BU*ۜ1��1
��r몖��u�=-��9�`�gY���s�B}?�"FSk�_Ψ���@*@H���,�1& �m#m-���St�4e�!���s���|�t_�Ff�}�(R����0��E��FE7�C������+�-�A3 
��%W��`�������{ުYrF���i'�$Y(��J��L ��Q��v(ϴ��*���v����<}I�+��~&f�����T��������:5���6�����G��=����b�O(v�x��4!�6Z�@��L���z�K��C�&72ʦ��|P����o�id�sd*�ۡ1e��*X�(�G�-�P��i�x6	,%��=m 3��  ��y�x��PSB�*&ӕ�bqJ������5E��d�撷	��e1ѥ��s�LA#㞣Σ��Js!N�	J8�ȧ,)��ɫ�q���3���jK$�BP^���	�Ė��r�Z4���h����{ݨGm�,"1I���=�4M���<�
 Z�sBH����zαY\��v�_!]�e����6�_��=�\���7�Z�Ǻk�W�x/�\�JT�=�"�}�ED1��%N�p��w�����;�z�
�!�ծY�|k7|V��T�:� ��3����ӶL�ߟ��/>Y��)K��|�6 ���V����GU�5�\+i��=!��;�]$^z��|�h��&����י���kw��j��@���NfCu�t="O?��@�������[]�d�;�e��1Њ�%�t~̊�����x�9;y�@��j�^�G�g���o?4䖌�@i��ubs�^k�ycs�(����:�-Ġ��ɉ��T��U<�k��
y�xl�l
����5�r�j�-�+	KD�ґ�~v�O�+.6�Y��S�Nw��xgnA�c"_��4zH�U�"�U㎶��[��JCm�HM2�2>�u��|���m�b������9yb/�Z����k"y�t��?e����;���j����k��E��G'ԛ�<SO�����߳ ?_vs�ra8}ލ_�0h��f�Z�/h��o����a�^kmN�:��Ys�U�e$E��co��w3k�O���M�\�+��V�̉��9-�:���Y���n%9�R�&ӥ���lw̮0l=$"uwOG��&��4���JE�ǡ�Vj������p�b���RKm5~}���QP�j���n&��v҂�;�m<Dx2�O���R�5`���N�GK5�w� ��3�p��g��1T&w�y�&�|fm%�����}Q����J��j����d�=֦3AD2Hl�>H���܉˶�4U%�����(�E"
u��5gZ��o�N1Q6t��9�p@�2X�L�[�Xo���=�)�#����;(Mİ�ȿ,�("Iְm��H�	s7z���Aɹs���J��~҂�c�F�BnFV�&���cD$�0���w79R���܎d�
s�)�UFT�����79�w>Bd�����LM�U� 	�^�Ynn���`�����<�MV5a�{��i�f/�E"~����-5�g�����x�rF�v.2���\V��ea�$��;�R'�ԩ]��<ǈy\����!l��r�R���Gn�W��{���l�Z�}����;��6����d���qv�#*~�����y���ڵ
ÌO�5�n3�Ga��N��+k��Y ���K���	O�N1�U~:��wl�as{4_�[y�eݩ;;�Y<W:��;���ؕB��ͬh�:�!�D�l&g=9�O��W:�Efʥ�t��^a��\����t���K��i:��٠�n�6�f�M��4_y��Q ���jX��yI��J���W`#���@�&�ƕ��^��u*�b���$m˓�GgU�3n��]dJ1���P9�a�)WQiy�˃7�L�� F,.�x��k�a��+��\�kS;��r���*7���9��>9$��%��i�g��P����a`�ţ�!6�T:�t�'�R��A�@�"�[���q�Dh�-5�]fg�<a�rڊ֮U�tpQ���~�e�Ճ<����+��,;��@w�>�B��Q�$/N�Rbwܓ{�������B ����ۦ gt�W�:�^�齧�����^� �V����1��nճ�vf�PNt �Yܚ��`iGw�ؼ�]l�Ƞ�{�>q�r2P���3�ׯ"Hu�/F�1���w��%/�f�[��U�Ig����qfxheb�j�E�O`�K�0�f�0Nu�U�?17�{���$\C���5A��e�8P����"���VFDo�'{�0�g3�LZC���0Q���8,!=����)l��a��\!:�d�m�h	!��{yg���L���ώ2�������7Wl�b�0�o>@P�]��,=I�1����-���Kh��>��Ɖ���*������V�pb)"�]z��ei��rl�>�x#e�Ûq,�y��`[�M�F�h�{�q>9x�֊��� ��� 2�����TF?A�s����e���]�G��,��\�SJ�E0џ�kf���P? �
��Y���O��US"v|P��i:vuf]�G#���,R�-�b�#/�O?�n$������s�y���)O����Q5~u��� �6
ˮ�Q��Ols�璉j2�� �tƞgiբ[��oi��^ ��n�� v�&vQ_���9Et]�J�E���`6}�0i��4i�0矾����5��6*�Ս���z��Q�lϡV�=��~) ���;&}�FP� y�*(�W�i�l+���0#R��F�����!�4�/��Y�K���[�U�xĲ7 {@R/���V�3:���0kh�zZf4���3.r�{�𠜣��c)�1�ҷ^�<܀�w���
+�A�}�sL�Ɖ�"�~�G��C��P��ci�����/�8㰟R�۝m���C^h�E�k4B9����^������kl!��H��ٓ[��B���|'T9v�_�#��U�Zm�
�P�x��:�1���ߔ�'�zd�`A}��]n�s7΁�"Ot���F~M!��t�;����*_7� ��JY&zR\����㳹1):2 	B�`tf�1��g5��wA�]��=`@��x|Թ[�\;��f�S�n<A/�&%��8�J^W^���-x�@B�P7�j�}�!f��qfS��P�,�IAcb��`��t��N�YT�����>a�AAT�k��]�dG"��(�s�}��g ��2d2Я���-g{��S��!o��$"~\t�Z9}~v��b��AQHr[{�"3ԛ2�,b�T&Ƣ�:�Oi)E�Q����*���ǕUp