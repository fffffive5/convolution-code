��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�H<�Bika�� ᬏ�?�{�M���t������y'	֣P����ϣs2�]�4 ~
�e�4�ߌ?�ҥ��QH�4�S.G��Ym�l�Teޤ�NJ|K9�|w��@z����]Ǩ���k�$�Pd�j�B<��r>�w�MM�G����f�K��u�"v
�;����'�ji&dֺ	�9k��Z_��1$av'��ob��g���U�[
����9!-Q��d?�ed,��WDM�R�r���P��hh��}N�6UFʗ�Dp�� ���á���,|�~k,/��
��W�	�]���Y4M�_�. T�E���Ř��0('�=�T�;x<�vtE�c�>��]lԊ�Y
�S��׭Y�4"�H��g��Y�a���i�[E����K�L�9�0�y[<�GR�s�U���!��4
%=3���k�Eb�`��LQ�S���mK�syP5&�c��	V2�D���3��2^$wr�z�4�Ʃ��A�f^�ז)����"��{eGonL*�ゐ	�%�d���.��`�l��e��>��X�)H��{��a�e�X[�Ȑ��[/��~ù"�.��?��i	�{����C\t�(��F9��PǏQ
�]ȑ�����O�8��0K�,-_���Ͷ7��c��R�QY� \I|�L�$$�4:��+AiM�ǽ���Hݼ���t?W9�JlE�Wzc��hO�諷!-���	ş�G���U2�P;��f��{�㎄x@w��30S,S4 �
βʲ{�UCJw�`w�Jظ���7���޼w���f�����#.ʄ��AP�5ФC�4��a욪+ _���dBZz��ח�o��~�e�pK�E}���.�f1n�jp����9��y�Ǹ��kg����_�/k}w@��f���y:�%`��B&,p(��^kD��E�C`����2@��X�=a5�x��m�e�o�9~��N;�0甗<�4R�����������dJ��)���]��EQ:J�5�*�ϴ� �����8��"�������,&�D�ir,���Fڽ�#{����i8׽����uM9>[ �4�U��;�I�� E�ǰ?@w������ƹ:��1qR37Q�X� �Q�u�<!3;�rI��v�NZ,������m�XF]�ǃ{lZ���޺�8��G�_�i�.�S����&)|�s)@�h��b-u}Jn.�'�2��փ/���.e-�m����r�ÔG�:7��>�� �_�,k�9���l��v�rX���K�����G��-R��;`l��b���u|<Q����lҲ�}�6[#�/�����1% ����flfpO�۹��!n�ļ<ɱ�ڼi�4?g>�"�cfI
&�z϶����ýwY��}�4�t?C�Ȑ��|9@�N�F��aZg6�x�V�A�| m2�
� ������ �0�4 ���CV��ūi�Z���	vGi�9�Zck�@�<H�.�x/|�M�Pa ��8���L��"��R� ��O��Ð�'a�ۀ�c�UD���V�aɿT\B����Ú����TY�f��<�Jֵ�������
Sg��p%�1%�8�B�
qt��J�s����	@�dzL�}�����rJ��14�[Y<�5�|¸���������ُ �;�ð��=�:�E�&W�:���`Z^�U#=��2��^�O�P>m����F�S	,��8;4Z��X{�Z7�@����� �M�JVF��,�����_�v���qx����gAQ�C528�c5w_d���]�$����X��Q�m�����p�r��q�;�����hG�a�ǻnS�F�&���ܔ0Ա��i��8xl9d����\���s�4c���&����'�u����1s�@Lh�4��)x��b�ht�9N1�+5�T���J�f!n��3��d�m��+8k�I��e3��� 2��8�܏���@9�Phka̟'6�(���]*I���j�[�� ,ɂ�H"��
�NMy��f�bjZ��"L�����=/��M����&.��f^���c�a9�]>,�6�z@,3�����&T x��Bf�ԅ΅�g»�"z3�}�B\,�������ף�9I��%�c�`�/��>�u��y��ڂ�##���_1�r���5$t��*._��s���Ȁ�����WN��	����N�r��ŗ�c`23�Jz >�0	��k�����Ů��zhQ7�@�
���ڜm�[�[�Քf�~�����KZj��� -#F:_�:�wtk܂3H�	hoy(e?����|��E��9�ĥ�G�+i�i��֪��^j�0y ��:)�������a�~2
c+M�6ZחD_;��zQ0��I�ϩ��B�.f����YJ��FM��8����̑�fUW��XC�ژ�a~a���}K$"����լ	zLrw���,p��4�|S���ç�ւCK��f6l�Ł[�~���*�n���_��~�*Y~&�)i���w�`�hM�5����}F�OJ<yʦ�������^Gu��l�~��SZʑ������Sn�$w�x��h��7|�̻� u��Ɂ0iiu��5ek'v����~���jU��>�4{N�w���5?@�Q��,��ƶ3�?��8���$����<Qr��z�i��X��`��mM�'K�)	�iU�D�?&�%?�_i'�D�4����Y��\
�d��o��g9�
�#-i��[���]�l��,l�`8+\���/e�r��pc���%jKW��k���.0�u� ��������DFއ�{��g�#1��D��3��}!��Y��xA'�t&'C�
.�;�R�`�Zo��M�h/��wUd�:��!ʣC j���
�
�l�_`?��^|x��_�sp��$�S�e���e�R�q(c��O�j�,����[Z�smQ�[�%f�/�\�#;	�~�`T3)��L�E�m����c��#Y42��WY���9�mQ�I��X��� ��J0O�Q�<�PN&��$�j�a�ϸ�ʛwnp���2��`�0�0?�N��PQi5,"��.aҪ$r:�+T}�g�}1���G�1�R�
�7�z���)Y<����!�Y7\}���$6ڢ�n�g<�%�D�Ժ�U�l�"(�|���L���ܹ���b�w,�������fg���C�)eg�u*0H��
�Tr���<���{���G�������4�<��6l��6��@��S��|7ԙ`�f{)���b^SN�� �s�V�Wk�.;K��>����e�u�(�s�:k�#�R��m{��2.B�cʬu��K�bE6��hj��^�
E�ӛ�����z���]��3�ar�����z�(���@c��Ӂ��g���gL���˳thb�p����2┹��(��/�J��X{��e_g�ߏdX�;���w-Ŏ�i�N"����-VX"8����d=8��IBVJ-������=6�ch5���љK��}����~ү�
�~� �_7�
�k�/	O�wI]{^�3D�j����@���m~U��64C��f���~�3���awTS�,A��!�2 g0oKK��H�a߮���;��E�|��B��O�X	N��"�D�y
�խ�o�J�m�bT l0T�3d��u�n�������Dt��R�`�4�[�_�w�r:hK7&��rbd�@���K��;Gg���9 0OA��&�ɠ��S|螢�Cr>rH��2>[:��'�SW���N�6���l���.��c[��z���:�= 4Q�%%R�Q�Z��DOd2��;o)��s=UO�B��c��i�q`��/��L!��5�E��Q��O�f_�u��r�k���`c�*���	�����22��}�ܺ�.J�������c�~Kݕ/H1��X����m�1bd�8��m�F�	{��%�f����о��>R���ȶ�>�K�C��Y��<�����ό	EX��^��RQf��A�.b�Y"� NS𖲷����>��v�F��NG�:n�"
줡�@�N5��~˺�vƛ�¯�I����;�hJG�%�<��I�@���j9�`K��OƱ &S�JC�G\;�+���Ƭ���h۬e��K�E�eH��$l�bJRcp
C$Fê�2���2Ϭu�$
b�}�I�Z�R@8��h�I�ึ-Fh �_��
���t�D�'"����H�������O�����ANa�! e���r�f��E��!��� ����g�Q!>�g��"��t]�9��ď��ܓ�)3��;��>��m�W�y�\è|7峜}-��<�u`I�>�
�hl{G����P��u�>O���F�[�/��i���wx�d�Q����{��&�^�Y�	��&�r��W^�nN�+��b�@h�*o�eP��n�Q#��R�~ϷJ�CЃ��\�ݟ����;��:T�z%�Ʈ����Î�^]ge�Rxl�X�?�M�
)c��	��U��U��eH��^*f�ӵ2s���ڗ_ ��.�o��}�9��2D��3�/_\�{�=�2z���|�b�d���}��D�͂�[�ls�в"�y�C�SX\��|�����S�s��g����KF�q
����%YG6��I��)`L۷�\�G�{��u[K� b|�|O���x�?��,\@���Yayn��1N�`j�1�Xpm��~o��x�;����a9cdv5-��at���-;��z�� UUQ*n�?�߇���ib\z�����5a/����_�l˔�wA��_�*�PG��n�:���_e�R��ĸ��_��Ӑ~)�˖�>fd��-��9.NQ�����O��!J�����"�
�E�f�Y�O��x ����3:{܉���3!��*�4s���eJ5�����wԂ�UpM?F�4������hb�3��P(ҍa1��*�7��r��
�v�6|�����&�p��f�fyP�(%�B�d���_��4.pޑ�M߿k�>�n1���Gvq���!uQ�n�XW�y._���_����*���x��cm�g��_���_���m�-j[������|$0��5�Ol��4���� "Zz�KDF�o�-+鄜�ţ�K�3=�����������uW��t�:zY���kA"um݁����Jw�w�����#�L������(+n�q�n��)�i5����)!�����Όι�WO�	}b�^�1�j�CW��d��U����ˊu�4C�/}�m��r-���u��,�Z�0���J��)&���NV-(������!{����r<l2M�>b''D�r�ƺ�0��~��k�@&�O.U�f�;B\��^��B�D��mB���HJ���ɞ�vmb�s)�1:�Z��ԉf�]./k"�ϗ"���4V'�~�,7�M���k��vm�L~�f��= 8p���z��v�Xza���H���Ӡ���[��y�b���qд\�GM �B��ϮpQz��ih�a�ʤ_�����ѣ�������|�2(�Z)�\Tt�%��J����:��P�I�	r�~LH	�Y���Ay6��,���o�o�>È�yB9x�� �)>��xXk �v�^���f<Ͳ2����5��.(:s��c���J���3��� >#E����M���#��n�M����T��T�c&�%0o�<� ��l��l�	�G�R<�N�7�,�14be��Ga��XB�-�t��3+��;��ŰR��
��c?x}�>t�`v8�2�u�2��f���q'5$�>���,Ls���S�<%� :�R|Ћ�?�a�����{�z�K��*[�is��� W{��E��2P�1A$��KvmVw%�mx��_��kn�)�S��������
&�($�C:�`�S�ϱ��
fi���Bѽ��@!�%	/[b��P+e� �1z6�c NV��!)��}�Gl��J����c�w����Ǎ���@ c��A�}�+j�ZлL��Ǚ'�m{�d:��u)��Zo�GlO%�b,��pk?� f�iq��g�#��k��8��E���y�ɐ.TIf��0p���'�Gc��g�d~�
��Ô�&��,<d-#c�֧o�J*:,�W!�4`��<��@ 6��r�iz֠��m��tB��1Ș[�/=m@��?��k��F�Ի��G�ns���Ѱ��a���ϥ*A����X8���FZ����D"l��y�po]d!ü��ݒ����S�Nu��'��x)�-�ަ������U�|��K�pǹ�C���5�dF��Uxt1d|�0Ӣʟ ��B��+�[~+V���U���n���\�1��Ԏ�O��N0�K0�~ay0�8��Z�-8���d O��E�����_�59��G4��G^!
?��h�!����t�qEC��#�6������t���Pļ��Y��#�N�h�l��%nѤ���ppߩ�w��7���ͪ���\0BX
V���*�Q4Ѭ�Tz���Z�F�94�����W�DLG�{1��ckN؅ъ~�bS็�+��t��Ë��0q�Dڝ26j�l��+��v���Iᯔ��~�ΰ���k���͍}��EV-�,�����:�-26]��nD1\�;H�nC\'X@����3���~�Z�z�����(���S����.��̵����W) �R�b���C%��]���,].�#G?���u�ɹ$<�Nn��#F�c���F�+��w������b�˱Nt i�L|�7���7jӋ���Ӻje�a����,T��[������h�b���W�a��N�]B��_t�[T�&�v(�;�>�Qi!Ⱦ����5�)�tR�Ǘ(2-h
uh��[���Rn6~;�,��?���KyG��E�כz����\}/5�l���7�j��㬊�~Ң�^�����ye����� [R�E�� �bG�ZY�g�hqGY�l����hK�Ǣ6�����c�to'�;�uT[��y�pTgW�Z��7��@�i!��s�u���P×W�K܊�?Oo�\n�Р�v$(�v�aH'�X}p
��BQ=�e���8D�a�+�����)2�/����8���j�r��	�̝Ջbmީ���s��tz߫�q��R�q(��Y(�F���W���.�blQ��cLQ��j?�y�9�c�+ȼ�+z �����Ø��`��dҒ�q��4����@�m�}CaS���#����k�}E���+�PG�k�C��������M���t�"c�"��kJL�T������9��^yf�+��>�mQ��	O��lr��
Td�Ը<wX�<rWk���Rs��:<�*���:���Y��a���s5n���S`#<o͏�³5�t�������7��bbfj��nF#E���(R�sa|�Hg�����H���ݵ =]��.&6-�!A�}��|��ԣ�\@i���)3D�W0��˕�v��c[q�Q��j�B�c���Z]��/�qҷ�_�Mt���"d�1�0 ��۷;b �M��`c�~ �.ٮ�r��oL��^/��9z�o���a��h��r� ��!g��a*���#Zm�{r)�α��j;�< ł�绠L��g4�6J��I���4O,U$��ΙY��~8N�w�BI}��$�~�1����W !�#&V�J�>�B��E̚�RG{�S�rX<:c���X�@���,��a֨]�~tZ�8�n��d���ڿ�p��3�:��%�	<�'?����t�dl�t�.�Do����yg�K���	7{ki_mC����5���ހ��i��ќ�:��G)Xjtn��H'���c�(�j/���{���a�y��ū�"�ks��]o�R
 �mH��"��d��� =��
Kb4�d]�C�b+�
r�p8��Ė�\鱹k�k]���I� +'W�*����ݺO��?J��q;���W	�>aR����V!����i�ٶ(8F6����`�/�K� �|S"�^_GpI��z��~��=���D#ڽM��A�J�W�|ps	.m��M��#RBO��@����%r������Ψ��-�>��ҁ��6>�#L�Tm�[�������P	�!yR�z�K7��cѿV�+�0�#��4�E��P<{�щ4	�]�]�r� �v�"���4�GN�.f�T�u�`���| yE��$мot�3�y�0���5ȗ����B�*Z�L�dM����P[?qs�p�ýu��6/#�h��aF��[��B��[����BD�w)/����Wf�T��#g�N�`so$fR~_r2�/O$�1�y��\R@T�/pjwc�Ck� S��[��!��A���)��#�Z�4X���G��Ɗ��p�;�R�­"�ݱxC��iN����#ݗ�Z��s�ݔ8�{�n�7-5����re�%5��!��_+�Ԃ�~#�}՘���n�'˔�/&Ҩ�2a��#��r�H�A"v#}�S���[�^O�v����y<��Jj�S�֬��R�8_׹��=���2{1ײ և^�� �����\n` {o���^�UVKm�@��^f��CZ���k����z|i�l6 n�*��}I]��3���';�����i���6㈶o���	�*����-�r��DzC82�(I2��aQ��E��%m����$�L�"�e�W��ˤ�-�5��)�7F%g+��!������{Bt�y�loz�b��+fљ���	��� �-m١Q\�f���]W\9X�1k��O.���P�	JD��*��'n�9��v�b�X,�����A�����a>?#��p_�ھ�9�Cca�TJ�4=����52����aŬ��BL0�EQ�H�7��@c�X,QO���L�l��b
�L�e��Y/�2��!gW(���9�	�����u��p����q�[+�0��}�A�N�R��K�o*N��,�~c���J�۳A��1c�_����Vjg[�,}���B�s��45p>���HWbm�Ȝ�&�"������ņ�N��3�[�T!l�Ǫ��U2^��XG���| 1S��>-��oK�\s�����~UһkZ5�a��\�?O�T���O���8%R���Čt�q��"a��m���=��;�}��=V��������w���l@��C���Ul���L��A7�l`9�iL Kyhj���d}�Dd�j�H�%ʁ�Ȑp��6�q1�[l�6���i֧�"�֋�N�j%���ZBHZ����N�Si;l��m�=dBE��c�ͥ�O���0�N�緁d���T�MG�;���+dˌ���|?~#0鐒	��J/O����Φ�����:�+���f b8M@��M����b̗�S$�A8P���bh�·��K\Dɥn��Za ��<�On�h������;:�@�3t*q U��7�� 	В�b�V��n���q8>��Y�yԭNa�6S�	����R�U#�������j]����\D%"���͍`���dY�ݩ�z��K�>i�f�����%��7e��ڂ���٦l���eE�%�ڿ\�������A�����y	�R~�����*]� ��ejc\Q�/èQv�����F'U�.]֩7�=�_:zHV�^�,Juw�B�
h�"򒟐�[���Ő���or
)�d���Pr�f�ә��t� !/��N.�ډm
ݨ`H�Wd-w����b�z	�q�(T%��P+2��Gt�,У�hӆ)g�p�K�<cB7%b��X@�Cq���J-��U23�U ��;u����y���������|��e3���c�)�9����
���f�Z�XG]ՙ�*(G�j}L�w�L+��K���IMS?��lu�Щ��氨� ���qս�ןE�h�4$DD��s�f�����	�~�
݉�� �v�����;(�sq��ⴒ���??ߩ�r">mHNy�%kb����띉����4�����4@��)[�Hú��$��{��;I<�����Ĺ|���n;V��~�*ͅ<�1,�[�8N���xFx��!,K����R�?��2�y(^�=����P���Nc��1�>@V{�o}(�#��f�z(�5�P2����ۑ	��ԋ���LM4(\B�������)>�%��qƬ��ny�:������X-@U;&� C��ӌ�u^7 \���C����N��I�'��S�2�p�g>�ڻ��U���y�ɞ�4>�#F�*���7��v�Q�jK�1�HA�<�W��ZR^�W�RKѱ���ԙ�ↅL��Д�C�͹�3�b0W��/��C9�v>���o���P���-�˶-���&��v�ؼ��ׁ�C�ʱ؊1�yN��i�cb�^�[����;L;���������O����B~��0Ciud��)���"W������Au[򋝤_5|jyV-H2�+!���iiOR�yC3�KX�Д*�f�xQ���o�|��!�]/�M�Z�kJ�(�'��ιa�*(6P選ͥ�Ga+;4�,3�~��"a��G�sB9�D��E5Kɢ�����}n{�>Yg8�Ѻ��D3CBۦ��O�<ބn^���o�2��3����t���aXr���W�4�!��	a;�}CO�kq���m7sCE�\��
�8�.�$�@zg�'������S�e�x��!Vv�"�⼩���p����� �XKe����69��E�>�s���Kti���)@��d��ܙ�p�X�e��t�R;�^�o���`T���u�Y�ƀ�yT����p�4������q��C^f/7D57�$�w_/Q߿�<1� �ذؑ2��kD�"sT��fjb8���󢟹� ���Z�g��8%3� {�V8�8f�,vƚ1�Y�jPt^���!�p@e�'��P*W��Le�O�R����>����$�U0�`cJ��{�8���O8�&z��En�2��O�X����S'��(AeC,a�#���|x�Հ�ȁ}�e]��)XL���%F=�������ͤ�ʓ�I}�_��h�`�)�Hu�̘A�gT
����ʦ��1�^�;��.�*��ԛS˞~��E�Հ[MK��g��̈1�-wb�蛡at�X���6"Bc�sCh�L=�9AJ>�y7��J��]�n;dc�����S@���`� G���)7f��R'��+���� <5�S��J���\��
�q|�t�D롋�z����;�e�7����ً3J��\/�������=���Ir6dv�}!Qԯw��,�{D��\!.-4�Y쐕j��Ua��L`�t��T~xVg1W�����9�>�ZaE$a�	�얕�ג䥌A���\D�ESH���&�QkH� $�)kq�� _B�������G�]���z�8#�Ĥ����|�j�N�n�u:r�QCv���[��۽��e_%:,��Oi�s h�ӯ��Q �nG�f����l��7����b�lO�����L�	�x�=��?d0�v"�8S�qg �A�\ܫ �_���jĀ�]?�^�1�yy݄,�~�WГhV�Ȣ�}�FÊS�����+#���H�e�Pr��!;������i��3]�%8%��7�l�Z��J��ɀE��M�>=m)9!V��W��0�����	���<��9�.#�"�Ҍ|���A�l��)O9�X^��h�����F�<C�_��������M[`Y���=�i$���D^�?��<�f_���ɛ�b��L����5O�VQ�%9�����<lU�t�Z����bp�.~v�&�-Hpt˝� ��%Td[�)9	�m�_Ι�Γ֒���f��^��hN����b�6��8��푠Ӷ�q�-�YpEB�n��г�V����|B�Q¥unЛ7n��V�It��ڕN�+7���`,}��bڰ�?0�������}�d��v��?�s$��A�|tәEZ�6�h,��n��>ܣ��g�gk��,�$Z�+A�� ��4��kٓy�8����$E4��/�Iy*x�<|�p>QT��Wjj�[W"ɺd��ǵ褂�w�|��>�8�-bdo$�����/��Z������u͛v籚�3�Rer���\�qG q�Y�W��{§�LI�%T)-6$���f<��J�&#x^Q����_y�/_�0�K���eY�m��nÕ���I<o��㜍��Wv�hΘ�X��A��GV|�n�M�����d�9�oAY�����j� �s0F�d�|m���w���Ma���#�s���F�r�B�m�����"e�*k�s��@�<T�H�槝V�H��N+�sV�k�J% ���9P��1kv��D�2���o��Wc�W0>g��yR�$�疏�Ȩ9���/�)N��e��B�:}�I*¼�������Ft(/eQZ�� ���~�g��bd�M�����L��Xm�����L"t03m�Hi���Q�&��F��ڔ\}\�y�AI����_�߸��4q����.q�l&@�%i���g���3d	e6Z�^�,I�r92[�	���#�BXR|E�����"�� |��p�N�g�Mc)�ipkq��KM�g��Uoo��<ΤQ '<#�*2_A_��v@v�x�=��Y�sWp-���h S `)��ߦ������˕+_�p���
j�n��V�~�څ$�j��+�A'e�Xs6Sw����\~+��]�#O�y�I��)B ��D� ��4�?��JV7���ʆd���&�h�hߡ3eE����(����'�(�
�Ϫ�4�0��UȜ?��q�F3�oX᧳j��@_�L �m|�7��by���t(����*I�o^�5�`0$��sZQ^ʄ��mNx[��c[62��Z���$@��c2?��d�!�d����v|q�S9��a��ew�v��������5�a�ӆ�݈S�dMt�K�����L���HxŜY�_��v�t���\ڣ��xf)%�	�7���B[^�H,�R��/�PMR�o��X��f&�V�W*S��N��tH�#l`ԟ� �l���lӓ
��KSڦJ;�ʶ�%7GE�s�k�^����e�t�Èf�a �Z�X����=�_ВO�%�S�C�3�)�f���
v_��n8.i
���%�3<pWE��/MU�3�WT��1�I�72��*"&K�4��xG���Hd_S�#��dN-�i���'7F�
7�B�qr�x}W$�����_����6�SI(�������~��Z-��Bv-:���	wz�C�r$V0�Whɉd��x�v��2��\����tS�W���'c��B����4�IGg5A�l)Ue�(������,Aѵ2�\���|��	P־rtx�5
�?�d�i���tV_�V�K�{�BC�m:U?Kt�=⼋��kW�������:6��F��|5��(�-�'��;�pq$�Ɛ�N����&]��p #��9��|�����d��5 �g��|T�hp�Z�/� ��9|Q`��LǶs�"3�tz�:xN1<��vn�$|��N�^@ِ����Z�0)xl
�T����;�V�@<�q��<1�����b�L��k|�ff=��1�
����$_���G���z�&�"�����Ruɀ�lb��	�I�ֆH�cT�@U�ԜI`'����P�<r#}�FE��:l�jI�� �X�8�BS�$0}j����S2x��wǛ�����\�>��[�|`���@�T ��䢗z<��@��+e�=̔h�\繇�[#�S��F�{�'c{rp�J���@j�&ㇴp��Ua�
Y��s���i}�4P�l��Y#d��#=跃��<J2���͆�É�
�m߆�=�R���$���ڱ6���l��sU	�|���$;�c��äbƎ؂ٚq#�r�z�s	��Fb`�ɀ�Y�ZK���_�:�/hV�Щ�\|�;UT��<H�b����H�:��JG��wO�([d��EQY#@�f�!4����5wqQ��9�u���Z��v��X�[֙˩���8�iKU���jҿI�1����O�c�
������ǰ�O��#H/�q�̮��%�E;q�8���Rn�J4�j0�-ǀ��2�eٺ��-��(�{�f炘��zm�r��a� ��Mi���t�$��` L���u�<�Y�K�8��ϓ�A「�K�����d���#���f�osgE��s�WJ$��#�U��E�#���y�1	J0�9��-�nr����;C���xb1��m��c� �'
����O�F�?�S���Mw�y�����@�f�:���{��W�d����r�`�V ��I�l#�6��g_b�{��0ц��D��6��l�_�5�?V}��"k-7������3�O���LZ�9峦����'p���ņ����/7��u����ȖkN2d8n|�\&�=5e�  �#g?:9vom��V�����,G9Xm5�Wʟ�Wj�]�q�y���s!D�_< �����q�V���m1�4��R�8O�:�
�L�X���صF�G��	�Ԋg̍��h��9�S���xn�GHf,����0O-F�w����P:�ǽ�b]fOƒ� 
U)M�����;,鑷	��\A ��8r�V����u� _E��NOk�g~]���g�Y`�/C�&kE~Wwx\���6��Y�ѴM8�sN��A��X.�.}���V$�K��1�g�QHU��<>TFe��t�Q��V���j��%ת��
zC,�J����<�}��s�x�J/�MCj���}��9��nixs19���ʒ.|{�y( .���_�E�Hs�A�d�R�M�z��c2��y��򡸩s�e)�v�ދiu�eͧ�^ߞ��(�����#ռ6o�p\у���vY�����T���m{�Bz����9"�I��fpN�8�|Z4`.w�L`e
EG�j�R�d��HA�����c�Y� ��*�j0���gZ@���M8��z��U{R�(^=T��W��)�Ǎ�a�$�;�Wa� bQ�DJ�:��%������;:ȥ1_���e�~?�QG\��Py��oq�R�3��=��7��SMU���B����i���5^��HXw��m~滪�C|��a�Z�
������e�5�b�yo^�S^�4	:y�c�������CZ���]-&��mtt�q����-����Y:9�E���X8���<�<j�81zc5��vt���;��u�l�#��9u���1�:D/�t�Hk47A��a��������Ƣ�?�ƣG��Guh�<	��䈧���5Ã�&�������� �?��U@����!�:�r�.�dߢ�����=��{�Ye�XE5�O_gL���? M�B��!�� o��;�W�,-i�Ս�X̐|redi�Τ�}���x�U��!�f��$m�-�܊Ne+���zd<q'0���>K�r��PO�OA���M�4d��2[����h�����-���b=�QW�3m4o�~����g_�J��'�oь��\+���$p��c
k��Hax�]X�l&��/*��N����!����0��1x�+��f��V}2�5�=��Y^�*<)����N~�BX)B��$P��m�w������Lk̋=�,|Ɉ��	��Ե���5L����jp߃��/� \;�O�?h�B��M�b΋��S>~�gt�����:i��<W�*�p��b�E������[j���3ZZj�tbz����֯<�?�VA�V�v��H����I�n�d��O`��]0���0�������*�꼈&��Ĉ���x	Ÿ��|UZ� �����#�6���t�n��*�HՀ΄�$��;�)&R$�D8B�b,٨ܰ"|�	Kl�R�i2 ��'u�q^�֧08�����z|(Z%���(����5�����R�I�/IU_lq�VY��Ql
�C|����˛{;���(0�<(!���x͚~�1�(6�G��]R��7tp=�aDV�I��_`+K�&hD\ja	�����4
���q�;2[���)`���Rz:D�t��9ě� i-�x�#��:;ӿZV�*
���H{��q&�d��9���E���.��%�V��!bh��~ZJ����XN��-_�
�k��䁡�f�N�Lj�o疃g�r�y�
|hC���da�ꄛ��-��6^].Yb�����H���I������n�G��ԟC$�%�\Ć��#�W%��k ����9rE���<A���`�ϾZ��6ͣ��j@��m���.q�U�������#��>�)����yB,��>�
��",�Lc�l3�(��}k��N��08*��N����hT ��j4d/�����%�c��'�b���e��RZ�wL���$��.�c�[��"1�LØ��W�}�`r�vG:n2:,�Q��}k�jF�고|�ޞT9-�rC�o3�^Lά�2�6���v���'}{�q�"R��P��m� �l~5��"5��Q��ǲI��$���O�v���>��Nz�f�L��^��n&�@�N�h�/e�0A�OІ8��Id���{�P<�'��Xh=�VW��9t�uO� zNeJ))��  ����y�n���!Va��>%m=pܶ�b��+"�qRk��l4�92��J���1,|��a������^b�SE��p]�XW����f�n��D�(���ڂ�އl�8Gs�뀫�Y:�V�^�ٳ��jsT­�ĉ3���0o
 j��,��g���ݏ`�I?�U��}i�u���ư��p"\(�,����xQ08��AMꭴ�o���5Q8�U��q��L"�3��d��^-�	/}|ӴU�B�S�#���M`�*`�jZ�I������G4OZ+�Ť���=���%?f>>�s�7�0E��/<a��aa6n��'���kL��coP�M�٫
@&�N�6�o�����5ٔ�)[ I���B�����*�f�7r%�{T��QH�:�y �mxjjNK���ړ����p��wh�u���_#��4�����#f�����?�i!��c��0�|�1������i�o�ZJx=R��~j�D�Dݸo�1ؐ��,�[퀻
��./ۜ���.ʘ�ps�������K S&�R�g��;�ύh56�49�Ss��֊:+�u2 �̅q�e�^-����c��/�;���ScJ$�٫7�s=䘹]$qwH3佢�N��� [����Y[���lh�UՎ�K2bJBsl�o)w2뛸���S�6%���;�?~Skr������,�|�;���g9�ӥ���U�u{Pco	��i�e�d9ʢ/����u�l+�.B��	Dy���r��d��^S��bH_�,P,bP���Ĉ���ٿ��Dl�W���	��T��*p�4E�����R���!u��l(*������IY��`vm8.�(���A�'��Ǥ� E��z$�4�V�)5/w��|���c��s�gCI��x9�2$ZRUz~� ]P�a�w��:>h�uʱ΢S�kV°$!�l"���ˁ�<�%��K,V%i&߃� A���e�K��Зi�s�1��{�Q�ِ�!.t�tko��?����G�;%$�Q�/:δr�p���A@��Z{�+'�'�pژ9W���f/S����YQDX����S��S�I�������^J�0������$jB�jzI�51v�I�K7��f ��#Tt�k���HT�r�ļ�R�b�l���|�$���j�H��
	��R|fp���eT��TJ��	>*LO?VXk�op4ĉ�B��d\��j��X��&���y��y�� 0��xc����`�{[�=[ww���s��
Q	hy�L�p�E���y!p�r%���dĹ�wl�::<���X��R���7IT�ǒ0�ࠞ�0f��QT`�����h�,{ ��7�W�K���I5�}=�����8ru��=������g�g���57��hc�T��tO�c��s��-��7��F'h�!���+X?��Ƭ�M/<�r{��������%��9E��_g���Y���f԰�o��4���cC��ZZ���S@�]��Z�e�w��?����u�#*��2������T��D�Igۧ�} �F{V��7���+85�0���N8�n"wc��7��e<����2z��ym�03��V �[�W4t�fl�X׏�Ŀp'���%���ۯD��:0�Ƒ,-�.C��F�-��S�"(���@�Y�uOac�:�lqE"x/T��+�[��\�ة��w�I�W��F������r�l�O��>���g��G�����(>� ��!��,����\��[ٳ�b�����>����.�5Sn�Lt��CUƒ�����ϗ	����ԙ5�vq��O&;d1'�m�9�"y-�������?�v�n����5ӟ=��P#�HQ�w��a��gA�@yW$Ŵ]J�@"-�Yӏ�?�����ׄ�t���4
����5u�eX���rS��L�l��
n/m&���)D���6��E�*��9�K���͖D{b]�
���Q������PQ�y�� �NM{|1��u��Ӝ@��>���$��~��p���x�r4�����9M��q�}��_b��}{������T��KpcE`j4����Gi77gؾ�(�����/�JD�'�W��La��t��I~_+��W"W~N`����6�o����uCD�6ëBni��Z�KmB��#��\�.���Ki�@�{�ZU�@�K��j@���Te�����2_iQR[b���i����3/�������P'Q�>R2�e<��flt�.e�8Nq�o�"�Y�E��r1���F4v�Y����fk�5��}�;ε��J�3�D@jz~��+�@ӌ��R_�~����l�#|���SJ;�F3\Q���/*��'�~t.p-���쐑M[���צ|�)�xY��������Zavq�@��(7`:R�ӏ���B���kA� �������I��Z��w֩+��ˀ&�X.,j�s�`�ww��=�z�0Ѱ6��$![��\�o�)ȧ�~&|\��{���hz=�ib�O{��v��A�;��i�m�=��z������گ,��l�,]Q|RP[_-N�+@�W-��4�yll�P����l�y>̝؏ Ō�b��G�m
�u�U~��h�X�]��~�1��Y,��+���pN+8��@T�d��7�e�qRX�����ީ�6��{�/@u��7�{���e��� ���B��)zѲ�� XZsw�B����E�b)���= �q�7�>px�8�核�-���3W��bӜp^��#�H�� ���}�M��6������A<l���/b�O�S}�[�w5E�$�Q��#i�ao��>_H� ������%a�(��s��0f;Tn�.�x��	ƾ'�a
0w⡙5��2-�Dd/� Lg�,�w��Y�R�?!'	�zR&�K\�) �EF:&cE����uP�,��SD���>B����;�9*�T��<���&��Ql�h��L�3�E-�m��I�X� �o���Q�l 4��ƄI���X4�buJ�z�)T0 /��)R���yt�h_[�J� ���6�]�}��:w-�>��Y�s�F�2�n�p�����>����	��-j����n*�f�s���Xda���㝏F�6#Ni�ѣ��jJ���3�������س =7��xr-7�-�=E��u3L�D�.���+K�Ή�	jR/�Y���Tf���y7�2L1�k{���Q2�o5م(4uG�ý�SI<Gn/���8�K[��;y�$V���Fg��_)��
��!���`�2î�LQ���A�<�HT�^�G��	i��{�Mf�����о�̿c�!$�N������U��KZ��Wm?��p�Skqy��73��3�WGNN���x�Y�T��)��ħ,���k��S��tc�д|V	s
�CK��(�J�H煺��v�(���ׅɤkE|���Z��F�5���Ne=d�΅�@������[�g�&x=��:����<c��?�PwL��~EM �:����}�k�^�����B'���'���ZA�=��E��Cm���G~��m�M���F,O��&���j<������csE�x)���1?Z�N��6��Z�|X�n���������V.5L�I�q4ԉ
�r�$|��dW�
%,�+��lA��[��;���ګ�J�͌����?�ƭ��.�ΧL3�i�1m�;-�`�e$Cq|�!���P�d����!�4 Op�Y�����XQY�	{y�q����n NӡGζ�y'��o:�.rީb9���ܸX�t�v8�i!m���Gv�m��f�y�ܡ�v��������� a��o7��Oϲ����V�0����z�H��5MkdԀ�e%i�k~��+�-L�ؒb��a�'������)C�Lq����{Ol<������Tـ�t�ſ%X۳b���"�hJ\wq&q��zs�,�|�RT�Vg���%<�C��&b�����U^9a�r�3TG0w�.��>�f�����hY�x�دoR��5Kr�@	��0>�o�2���J���|�bO=q�0�2�ҙ㗔�j$f.�~�ȁ��K� f!��Y����U�V��s/������  9"}P��Ј6;l��@Ʒ��LK��tK�[�X6��W3q��dh�e-�Ҝו�{��c�p5kw��/�;L�3l̷�D-������͐�Uʹ���}�~�5�@ �.8�o�_�Gn�kp	���4,�lh�*
4\j�.����j�|:��H*e{T˝D��F������\ܰ���?bک36����#\T��td�� E  ڼ^
�$orQ��J�|XY��رX�RR*���������_o�45\8j?�O2A�HԒk�=�Z<<�l�[�>�6�B�@���|�b�L�۴}ۊp]��R���6+y��7h�����wk���#����7�
��{!Cn��h�r.�����j���r\�B���ϔ�x��ź��7�*i.-u��s^v
f~Q��
��=T</��Rd8�̤�[f.�࢓��K���;B���T�a�
�x�ھ�sZHX�!��zb_�!7F3U������R���B}�9u�5�#'�ݝ\+�>��IzDW!+�X=�Ɍ�&�!0�����)�V�'́B>Vk�$(��	� �T���h׹��W���m`�	S���v����6���ز���ς��%�IOIb*b���(�(yU<�ƈ�P@��b���CE�Splh��?�SR
x[V�:�H��~#���ד3aR������Nb��Pݍ�]��tlJ����t��@��0A}���bW,'$��nm.�\G�>�|�`�����lcߖ2�HB4H��У��'���� �4��_4~�[�"��9��*A�d�����D/�Թ���W�Ww����W�*j���� dF��Բg�6u�&�|.dp�IL;��0O�����o��K��m}Y]{C!�R�AT�]���8�D��n�Jm)�h���t��^W�v{𐁯Z�B`�l,`H%��7�^������H'l�+Z���Uz9(�+��1G�	�40���^)�^(�gПXV��/k�8RI6>�����mH�x��3��z��k�]�ɨU���6�l�O���?t�AL�R`�g�O�]V���y�{���?٠��v���J�[ېt�Z�-dႶ����B�2��..����z`&�X�oD��	��@�\ ��U:d��Z.g���S�"f_y�{;��IV�i_��Q+ō@�+�#uNO��g�3�z
�XEenS)��}fz҉� +�H��A�\һY����`��Q��F�y�����Jy��,m���9_�]��I����/{�w?-��lP��T�qò��&59)ɝ�"i^�JAȧ�{��cW-��;&5�!�����Ô�~O���w��ձ~���Dw�A���4Wm��V/�u{����fa�`�t}[�����_��=�t\����ٱ�}�0����-?��&�~EO� b��&�Ye���)"WN1'V�B{�g�䨘XM�%L�`���E=����D)��Vc_nV�N(0 AJy`p���E��U������-�i���܁�)�V
$ܳ5PI���N-����R�m�Y'5�����l��2���X�EXXY��Y�f<m.�m{f�~�-�6P%T���R
-�x<�x���60+*�a0;`��.���`:���*���SY�R���Q����9���D��ֽ�&�L�lnb)h�5Ҳ7�P��~�f�OoB�e1�àK��<���Ed��\�Op��:��{�@S@�� �Z`�B�����kP��xk�c�����M�""��JlKnߙp6'L���P��p�!��AwM����'2ٜ�}LҦVG�=�����S�yV��E]91��9q�e8$)�������>�0I*_� )�Ԋt���� l��R�,�wxR���VqJ�c����u,� ���^Ó�Zn~���JH�;i�@g��tj덎�KO�*���$�S%��z3�W(������5�jd�v\-��r\8�~�	����`��<Zn��ע6�KD����\Owp?�u�rn�,B�U�w��V^\6�
|=�`Һ�꿛,��5�ߏ�@��/��g[ h,'-Y=b0)��|��g��":��Γi*�\�:��D��$
�	>x)}��;��0��o��������A�P�^�m�B}�t��qw�S?І����4\�I��%���\��3��}�Fu_�S5�@�U8���U�s��֌����%=������L����û���ց��.���7Ǻ4��
��^�����4d����Q(���ے>jG8)\�`�2�m��ɟN����SǄWc���h4��{R|N��b�A_K�FS�:K��jsܞ勵76�-������9:\Ih�>��������4{�}����`*ч	��0
>��6?6T�z8� �q,'�Or�g���vֻ.�=�Ơ�l�$����G���AX��Qc`���R��O���p��,��.-<���S��،��z�\7z$=�$R&-K2u��~}"c�#<��@E>C�g�'⑦����Ʃ�ܚ^���_�C1P�r,쭘�V1�~�*�b��^!�H��>�6v���`w��ć����B*4�YI���)r�"�)p;�L�j8��-��-4�{�&7�A��@�T�ǖ�d��xO�ۼ�f+�5n���KO�ߞ�=��"�zs�Q��RO__�ȱ�9�ۯt��`���D|7����?� �"0p�rh�q�)�i�����R��a�QS!�Զ�|{0�Вx�L�h�J�A���,,��xzS_`��u�@:B>)�6���^PB�X�O�8������l�U�r��f��KL�隕b�AC�]�ۣ�e�)�]��I\�/-;��Xyq�����5�,"��
�V��_�B%���_�����wW����ٍ�qA�����B7N��u >5} ��E�N:�u�v����m.�41|=u��T2,#�u
��1�9WӆQ�H"��yAE�e��l��6�g��-����50���{I`��h㯮%�(��������t�ތW���nΝA�z��5����p�Cʘ��b��K\�i�� y�(�pU��-1HAs��dSx��˳��:�Ք� Q	��TuA�~�Ű��K���5�R,Yg�h�\��D�������F��XN��i*��9h�޾EQ�ס��3y�o�?>N��~�ɔ�i��@�P#�z��1͛m���2H��'C�$i����nb��ݕ tg|��o��R�<�M7M�D��HG�}���S!��~�m��ɰ�R�
�u^&դ�j���"�(�~�M�t���"��6�0$ �,l
ݷ�M��HHϠ,tKO��`@�Y�%�"�_��#���Y��VSD'��,�d��\�{�eo�B�SH��ƀheA��lkyp���0���SV㿂%ۄԟŏ��Qf�R�Zb���-�l��+o5�N���"�� N	p.��g$Lp��:��� ����p��M�qh��Ne�,ET���F&�/�NwM���:����o�d�,�P��\=���g���	E~�)�~���b|]�{�G�DJ�!w�8�O>eXA����w�!�����ٰ���'�#�UO��B  U��\��W�vW�ɗ��82���a� �B�'�[1�e�>�Ԥ����/�[�i}�a��R�Yj噆Ĵ#&4F,��qH�;  ����2����!ܲ�%x�����X�����b�6�j��s1��9�Ա���G�r֋<LO�{�����'�Ax��%�>�d�_�M��L"����f�t�oݣ#��)��.Ù����)�
�ZC��d�n���Rc)���ƕ��N��J��)oT��.�D)����Gt햅�Y� ?���b��|�(K��d JG�`�1�|N:Y��u�bo��]ش0?��ݓ����S�'�6�d�	��0h���'W����ݍl^��;��z	K�c���s�O�5�p@r$b���!�����4��D���G6,))��]4�{#Zn�u�оtW���+J^fD�6����}|P�v>B��v�ť=�l��q])�C[�\��|
�UvŊ5G@��̘텷����M��ݨcna��q�)�n�./��k�E۩	��ؑ�A�/��;�ė
�j~�U���*B]O0�����GZSF_o6G�m<|zS���El(����	� Q�*Ʋ��-?�F]���	~�̘,�Q9տ'�!gm���ʡ����,��aV����	#�A���=�%���!˴rϼ�6�-8���ʥ2�	z+\�#�ރ�j��\�`�ާ���Jx��8�� �E	H_!M.���-�ݣ�/����֧0��U2&��X�j�[2���w9�r�X����J����)ñ�@R`{�7�[��T��U2�L�gT�s�0a?�xLD
�h��`��|��P��N����d�o-��9�B�5��3� � �ш��,X�!�km��Rгs�O]D�b��tvڨL��'��;���>���Au�������T�hn�o�8���Fg���,io���i>�P{KC��;�lHo������ژ��eלX�;�t�d�Af��n�Q��z/�����3��9�]�2��rs�2�}�n36r_��<��j���נ��!H%FO���a�.	7���ȗ�%�k�Y
�?�E����^5��>��O�
��;1��k%��|�8��H^����	!*�(Lf�mUGE=�6�
�u2d7f��?9"���������}� ~]3��߿�f��@�&9�.�r�f��-�:���J��{��'��zmG�0&��<!�{廽�
7��=���6�ޝ�Kd�i��~��gI����K�����/����_䰢�⾐-� C�׷`�'�&vg�.dwߪ���>^Y[$���;�+��O���ִ���+��}|�(��駨���m����b����'L7!��,�.G?>9�)�)�q�a��M?��\��p�v[C���̽���NFz; �=�J�|�����em�4���,�Gl=��m�ԅ�>Av����K�>�����i�F*� �� ~`y=(�\�2�rJϳ�����)��#�J9��I���u8����/Y�����!�]7���9KfMD�N�EZ+��ׄ:�3�6���|�Ja2SQ��n��(=(�J�!D�!�"��C�fHi�a��fa8)��)��Z�ǳW�` ��*�����,��0o^�;ׁF �n0A���i�`}H�)r�^P^��L ��u��z�u��O��Q/���H���Pc�}͢)����x�W.UosʙA�5�c�� .-(��W٫���s�����)/��*QZ&:�8���GC�H䣳�X��Pxs� +��a��6���5�+:`F�r�s�ϛ�Ii �m]�m%�B�:�%��O*�g�i������I�0��&{��HfNS���pKi���L1�.4��"Yo�Ց"%����{�	^Wo�@-��sN>@?�2l����Kƺ�3:�ApF��"����	�%���d��5K]���t�L,ϲ��>~�ɯ�j�8���=`Ã�r�Z��l��_�陉`�97�W�r1X	�(fb/7���鬓Q*m��Þ��d2���$ߪ�sT��و�_����3�_����^��=�9;9: z]��;��cq���>�*iQ�Ykw�"X�a߁�]af��� 8f�rF�������� ��l��ʮ����J�ra@��x,+� T�M	�!���Ui�6��v�VR�Zu3Ǔ�:���L{lnT:�	҇4X?�n_7rn��<|���w��<{ea��Y�V�q�����K}W��%Ĵ��1��X�H���]�M�K�{@���{��ʡk���H�X���w0D1���ľ�{ҕR��Ub	��:)c_�=��B��;���&�Z"so��{Kݖ�E��[���N���z�g&�u�?���2+@�0��99.��B@@�N�4U<
IJJ�`!��Y���k�_H\t	�R��>\)P9?g_(5�;�B�-�ʶ	��"��Tv\���r�^#u�S�uEb���T4r��2� �%����rMP�󈌦.�2����;̼�র�}�þ�b�D�
<v-���8�س�75��
Ҕ_k�M}�-/��$�Ŧ��̴�<�s�1���GÀצ��
���?jq8���6����K�Bg�]u��Td͜f�x�s��*�A�QplNm���m����Vh��:A*� c� {�G<��Bb8T{�rZ%i4�$%��c�t�w�*�9�o���_�Ǉi���,�|y{b�q:���=�'R!�Ds��q����}t!�l%��"��T��|�sH܂��3@�*kM�����5{eY�z��a�~�~NtX� �.�o�>h3=#6V�u��ТDt�]�.�cC6x��+��m��<@KT��@��Rx�Լ^ʄ�q�Te���V�IR����p\1�;�S;�hq|>VC���C����)��v��7\�x�se�q���$!Uڣ_*R�9�%���4\s���2xQd��'{�IG����Q@.g3��<��Nd��g��G�O1"\��h�KR�&��6u &q��8_f�Z����3�.�42��e�̓m�x_AB>��c82������Ieܿ<c�Z�+VA1�^�w��Ϟ~n��D~^�R�OiKҔ��#�R�8>���]�`�wԍ5@��GS5�����rh�eU�݆��L�=��y/��څ�_�$�LJL�9_̾�x�ߨ�#΋�S��rm�JαֻqG�ώ̃Hi�JGu^V����8�.��V�����i��J-���ī��y�Iu�ݩ|�s��(�Ed���S��N7
#Jݦ�������U���d��p&o�u���h.�2yY��c#�Qg�R0r�lȮD$<�v?��=���c2/,K��Bi3Ґ��9����)#����&����|6q�ԑY�$#�  �܊h��F���t�1!K�|}�vĳT��!�'�G2��Rm�g(G�8~]�+�$|C;
В���_t��a�v�K; ��P÷=8���_)(�[�HU�퐏x�ż�6�3���h<"Mf��ܽ�O:�4��~,��W�Z�5v�R���:�1�H<�ֹ�G����X�*�rjC��:�s���nja��.H��еv�z|� Wa�x�Z��Q��J�)��h� ��V���?gN|gb�� D>�l}�G�pA�	>/-��T8�-��Z�����"W�?'Z�re���T�:R"F���&(��<E��J�$�.[�]�B�J7�)>�_��S���0e �����Cr:�����B�n�2�'�~a;)z�$!��l�*�$�ۆ!"Ah!�^d�ۑm
hH�]�ݵ�� ���/���BRJC��}�[Y%2�;6�U�^no�B��:�����f2$5��2��!oy��g��ˈB�l��q���*��y�b�h��,�����B�; e9�+�������n�	��*�d�� U�3�#L�#0ҶD�1�r*M�bƆ��ߎ[P0�"��� (q�M�l��<�>�m�8��b�6#��f�i6e��U�;�\��1C$w8LڹF��>�4zd��Tl>?��#Yg����Y!2>@�� �OcE�i�wj�|�1n!����?����)����~r�o�E�'×NTFK�JW�dCǇ2�ވ��r0t����ȕ>|kn{����{Q{��0]�Y�˹M�q���%']����9��7M�B�`4�jU[�l^�%��
E8�����~�Km@�g"	����s���_[i��hT��\����8"������a���칠�`�Uh�;+JR�m��<����c�m�`��^R��O���
��@��gCl�I���3Q��-�2J� ^��̹����N�	Oϓ���<6���E�a۵�xS�N�J~����I��E�^E���F�p���5���N�bA����&u��8|@y�m�T!/����`�6��hS��F�,���VP�e�%N	:�΍�/FYu�6�˲��!�75���-q_���iw�!�Ù~���M]$� ��՟�92cL���+X.v{;px"���8iNr���?�+�N=�����ԼG\��[�s�����γX~�Ug��5Pʝ	��7?v��/�C���
��atwV�o��/��J�#�J�#z��n6/S6ahpPEh�P�B��\�YEz?j*h@�u�=����>��Zu�B)���~a�V�j����+�<����bHW[1Pg��#)��|'I����,�t+!h��ʚ�U�Ô����u���~����$�b��`�����~��k(�#Q����܍��+���*q�a̩��O?/-U��B��>�J�Za���:\oD�	м��_l3�Oeb$�͍,c3�N%��k�s�#���;�ai��h��$�j�u�X�;�y!��S5��B/��v=�E&]��z"�2d���xmG2#���e��|���B�ml|�[c�e�9������GN7���Bx.�͌�2x�N2ԡc�?\ueocEc�r��eˀ�J��cS�ߺ��y��]P���d�'^6o��u��~p�q�U��N��I�0�сV�4�*'�7��O��nR�n��,�9�0]`������Mt�5��V桷�N�1��A������oP���M�{�������Ձ?S�kگ��;�PY�'�*	���}4�w\��W��P��KirV�+���og��ߵ�>O!�6)��N�J,:\.��Sin�F>N���uӊۤ�Jx� *�R�⹚�0+K�wm��^��s�^~������߭�Ӌ軍$|c?U=Ĥ!~��`@�%�4��Ԗ.��L�9�⿣}Mx6<��E������1�Ę�~:�02j�9f�����`T�9Z�B��M�(�oe��D�M>��F�f�S���Y���z���.�'7裂��,!����6ݩ��$dz�V��6LСo]�mEM2�?"�W)�-��/��.�
�$���\'��a�▞l��ҳ�,+@��iy-�Cl~'��^
" �_�T�Ű���V�n���K =�k�S���ڈ6���$M{���)�������\�_o�����a��5A��3h�
�/EȈ��v�{�/ž��
�FG���������r�y�:Yع�dmU�b�����uP�����wkQ��ꤊ���� D7V�'��uHY�ge��g������B�i�h'�DQ�6٠e�G��#@&�Uq��s�ʸ�6� ���Y�eQ�h!1����C,Adam��:�x_m��3��Uh�9��5^U�E":G���i��)OWc��rr�E���Hf޵�'C���Q[`�HW�RXV��_M��o�g(�g�m}.
V.���V���~��y�L0Ϡ%$(���P�9�<�r4c�D�4��QSw�FY5#��M��b�ns{z3������|�FmTmF iR����pSa9p����l*�Fu���5�����u��*�����h]MF��^��h����ml��_�f�M�E���	��֑��kol�Wn�h#����N���%��n~cz���~=E�Б �ѭw���l���XBL$U�_���뎥׮nl5a�2�  ����T�
����K����Е��ړ@��9�V(��Ɩ����ۆ��H�c�/�Yhh���Gt�Q�T��v�ʰB1�v4����(7����f ��ǔ�,&Y�8����3��Z�i��*�bx�qn.l I53��eK�Y�_dSO��#�ĵ.����w�Fw�o�">�%�M��MDA��x.�����%���Ҏ|1�����E�j�%�o�!*�����K_�o����N'�v���Eٿ�2@=������������̰��'��B]�#r`eې��}���;�r�I�`&x��b�b��SK��:���T��	���ה��1��G���?q�'��s�|�����_���8�Ov<�=��UaԻU�5��ܨ\�7WP�k�`r�,�E\�/�[�P<�: �7q�_���<F�H��~@-��m�鈆�L�6Jz�/��	囮Q��4<��
*�_ �����a�]�#`{55�J���>L��DB�tr,��%Kz���x}B�*/ݻ=�sj�{W~0��-hq�vp��L�!���,�I�H9��n��=�pw�oFN鵻����ƾH@gM�xg�_}ca��T-!��G�m+��T_G���4��^�����z_N?�=�sP�|ƴ�]M/���t̀F�_�0�M�6�2l�1 q�L_�gtY�R4��=���P\σޮ峨�w��@��)���q[g'�P�:�a�K�]��r���b��'�P�t���ʕ[DjH���w�$Ti����.��s�ד��'�֓�������]�=qǷ��C9Og.�dR	"LNM�=�$���eZ�)�S��������, ؊���$,V�s��'��D{�$�g���"z`�VH�����#��K�fc�l�O�v�g�䧾�$^�F� ���n���+��a���K@�/�S�febu�F*��G7�e��l�p�m��Q��@���{�F��
�
%�g��R)�i�Z���[�J$�5Rق,�x&�JF/�A��c�ٮ�%��i�n��)��*@M�|��{�٩��x7�l�4�N9 �gQ5^K+[�I��P�s�>�o6-
�}���#��{�Ncݣ���"O�9����x�؞�Ӻ4�ľ��+���<J0E��AF�p4;G����ܥ�z���"��P	x����f<�L�����l$��-]����|�##�m@�&�)�i1��'�2����xZ)��re|H	о��̮XGh N.��#c�G�,`��Pq�1p���~e�]A��S�ё3}�w"����}���E0�S��G��l�aE�VxI����rؗ��l�L�tl��ɵ�g��\}A�!\�T�x#|�r'8���	��MwT���'�̟���Ji���`n��p��ڇ�NЀ��Hp<XF��VT�� ���i_4�2F4�xq��Tk{`cy
�nTZ\�`�#��qm��EVh��pbPwj�R��x��aM�8� �5�\`[�_ApK�������Ȉ��š-4^>L��67B�`���1@gK�.�5m����`ц�����ܷ�d{��w@F�.��3J׻��3�*=Dv���Å�-�0�8� ٱ���=~z"��Z߬�V���	�  ��(E�!BJZ��Y��3b]p�R�(�rz��I|�ۂE���_F[]<��~̩h�W�#F5�X��A/�b�t�ډ���6۩��K�->獝/�J"");��!O�s�y��s��Ġ;7қ
����~Fm�a`A6f����^���u�g�a�����I���2�����9<m�W���`"�1�}�@�4r�$�#��~�~��	��G����Li��)�Gf�WW�kƈ)��|^�\��[��p+1/Kת����w�Az�QWJ��%�A�2�͡�����U&F��MA� ӣ��᩷���:=]��<�94�Pk�J'����N����$��=�/�mE�u�3�9�/�D8]���~ܬ���b5�ƨn�й�RT��� #�fj*t�Y �s�_C��Xw=O��H�Ⱥs�{t١��rj�\�~9���{�<B+�У���������b'HP`�_+�7`b�hS�&@<�/$�Z�|�(u3�. �ق�����da�Sj2$V�0^1G�¦��L�j[ڒ�g!r�y�� �z�(� rǥ���Y��ҹd��R�8 ܐQ�pT=*u�yˀ�	N�w�e`�_|���QR�o�QOV��L����|�D k�f=��䵍=\#_�v�8��p�"d^���-�7��#�
���|ǚs�L7�o%�.�4��+��>+�\;����7����t�ec�+=�vD�L����iTd^ϥ�w��q'�^F%p ��3t��H��7�}�Sz�Ն���6@�㝧'f/��$@��5�ܐ�R��I�{?��0Ά+��hI�{�Sb��Ca$\CrVK��z��1_�X�`��AL��b:� �����AWx��?��N:�\(m��$%�Ύ��+~�����d~��L8ܸK\s�NR.#��G��hܢ������	���|�}~H��d�ց-��y�<����ӏ9���&���.t`�OYς1d<���c�2M�5%���MA����&L$i��L�_4Ѥ���ŕ*���yĀ=!�(Bk?�qx!co�6_�R��i{���*�u�c<J<Wk�s��G�%E�^�����yU�!�;Hw�ZI��B�U����<�J���n�s�m�$ �jՏ���◭{�t��MfAa�S�K�X�����.c��i��O�.��fI]I+���'�5{7�����P��� ,�PSC��'J�>�r�[>9	5P��ch�-�?ۭF�>�V,�".U��G��<��=�H��@���p���$Q|.k�:d�Q�N@mr	~'�����UX��[����2V���J���M��!#�3[�!��0z��hZ��Zo��p�*C#���fF�Κ9��E��-�U�A`��m1q
OC&l�"�~<�3&dmڧ��cU=��
+%�T࿫;[3Iw�"���GMpL6.����%rzk"�[�žc�t��e"�=H�e���Q�[�\|��G��l��>��YpfP��[R�(@(���z�z۳!׉z����hy�Xc�	�]�Qڹ�?��z=i
>��e"��ηJ>TD�3)t ���^[m�ɻ�C�Hۢ˭O�i�8��;Y�$Qy���ͯ��{W�+!�y�oD"��l�W�Ӷ�Ɨ�����$~�a¼I��	��̫ZE���sb)����±(=�v��K�&���4�c�+���wn��Z�hH�(Q�:�����"|��H*;����,�n~�X�k6 `�i��̻�8t�7�T��z��]g8���D�Q�^p��R���X��/un���|_�A�G�+�0v2>>@�F�m� �}p�TT���==�y�Q�]9z,��$�_�d=�E��՜w��rC��r� �_,�O���q�h��ܘ�cn���z�q�'su���\�*�}y��s���;�hN�V�Z��9�7�F�"�=.�P_��I˂���u啵����H%�3/�͍��?7��l��e�k�w^���`�nwb�t��y��agڹ�l	�]C��˙`��%3��7h���5�)M9�*2`���I��wӞ�p������qy@sQ��;Py�*$�R��}�f�mwi|�N*	��׺�(H݇��H�c:����h#	[�����ј�>S��'���-����^.j�{�'N�IZ�8�k	|�+��b���*�-����5h�Os_`0۾��b���Ǐ��`^�9���#Ѧ�M�A��;���. ����]�c�Ri��.Q��a� 1�;�=�;�p1roO�r�a�º�e�a.�c�N�(�Up�^�}��z�#Nr��&8�,z{�3��i%�>��3�#��fr"��(�WE�{��vi���TϝCݑb� Е=s���y�OE��׺gg�"D/�/C��"��#n�-!a+����j��)y�ň\��
�p� ��<X��3��b~���Y������1�Iwv�Fn�R3���^��S�4�
��fU	�G2J�a��1�O4�����Rd��֒�b���<�}����-���D�T�yp����'�9`յ�i�Y�&������	���[�����z��Ж�f֌<��6�x E�n<	�t?g���^���n��3��&{$	�Ω�]y�R���w���8um)5W�T�/~L[|�p2vQ%Щ_�4t�Y.㽗�h�֛�p#�:�Ȗ6���a�6w%����R� $�r�R�7���G�(��j�X$3p�盠�)��eu�1,uj��_� �'_N����؇����H2.��,��PoO�.�H�,��jaU� ӅP�x�PZ��=�`�y���{�dr�U���5�D�N�ac�s���{5�C8Ѫ�ѡ���G^�=�[��f�Ƒ ��O��;����0���eֈFT=wL����O��']SAM�7%�R:F�-k���{���W,���=?\s�c�P��Mβ�%�.r��I�`��N�F�X�ӭ���E���3v�B<
�GћDk���|�t�6�?�c?4?�t�֧��u�H��gaQ�\�~8ԯ�F�~u�"��� � ��_�I_Ɂж�" �ɱμ�u��Z��h��.ou3pVΧ��	aY��Me;T�&�����v�@�S��._S,6M0���O�9�
�d�u����pf��P+GN��X���7W3��i�v�_�����#lRd��&�+�_��1� ��~��H�fB�9��͔��8��{/>���7������ݠS"] j����`����X	�^i��V�j�_*���SE��ox>�Hg���N������CN'������eؘ`f��)[wC{??���h�<�������