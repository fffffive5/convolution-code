��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L����ʩv�*z�<�@������ ����*)��]K��lӥ�'D�a+�NABٸ�\�nyBt���t�x�!�A^TN�)]�
�2b�C���n'X܀�[5�L�d
/W?�9�:BӖ�
Q���pz��=#����)��H]��=ѝ��QJ��]�������l��* ���+wW�e0c5�	ƛ  �G3��U��xiv2���"�8���\�^2�;~�;���9E�*�7�d�m�1�٫N������]�y|�s�C贁D��Mo��,k>3�e�W ��L�����F��O*���=2)A:BF`ο��ܐ�(5*?���	�$IUc���;��|��#ݯ��_W��{��ۡ�v��Q�vg��g\�?)��&��z����2@F=�ފ�F>D�}�c��o�g<m)S���� YЁ�)�N&R1#*X)�1ټd|��^sh��M r�0�S�(�G%A�WB�4D�i����X㔗w8�~o+������U&�]���ꃲQ�z;{�2k'ʯ
`5Wd���%��QIRR!��'��~>�o"�wg)�^�4�_J$�Ԟb���lÜ�P�zw$��TY4dϾ���*�:��w���l8�l/ahO+E����	�4AgKI��1a��43)^t �W��{7P�]���x���&'aL�}*��zf�݄�P^\��Մ+3z��#��"ݑ:й�F]X����/U��a��.�9�*�4����[۸/������|�ݗ�(M
4-ɖ���N�)$tL���{�55Gk�Q7���4)M׊�0�Tk��gXq^�P_a�O�X}�*��G�Ѩ�`:l�1d+jJz�9�q�$]A���={�"��+�aÊ�^�+�1����ӂ���gV�i�� ��mF�c�>5��K���-zQ���a<�8��V3@�-B<��k3j�2S���]�	U�3�Ss����:�s�f�l�IwA��YZ*�xL������2+�L�i���FQT�р�{e���O� (plQ3	�A|X��ސT`6����
��nsԬr{��F�Z�K8��9�վc"7��~��q��e�6��� ��c�SDv�*qVΤU���,�G�֮���L�pe:���/<�6t�F�f���>�}�my�{����d��.�N�ݶ��_1������3Cߢ%ۨ i_����(��������B�����v�2vq�g�
zm4�C "?��f�b�w�R����|�]j�YS�
4� �s����SݾO�B_��;')Q"��y·�����y�C:��{`���q���*�Zt�`rE׭^�H�u����tG�ή�Ä�	����p���n�ЫRϣ��7�'�C����b�j8�;)x��?�����8�Q*[����ly@�ł@�ؑ�� íǫ��O1ܳD3���	����~E����,���0%g��V�ܗ�!o��z���b��[�`���Z\eG^���_�!ku�y2WID?$�iYa�
	7hs:6���y4/Ϙ��|�Z�P[��D��9���D���>�ۉ�"�L���g+��o��
�b�����Ђ��d�BNP�et"�|�LV�s&���;�����ۆ�d��j�w�T�_7��Ev�)ڣ��h�㦡�<c�YY�x���/6�{.q}�jT]I��/qt��qZ�����o'�*?�ET>D�Y`O�)���wO`e�Ob������4�"�pH�u��|F>8�3���Yh���rH�V��\��2�ǧ��L#cc?��LOVsn�.��X��8o�`���1�pT���9��L�4�������q��D�I�<f"��'�u2Y֭UM�BX��D���ɳ-�@�t��M�4	{��\]q��7xa�fyO��31{��N���o��eE�-��\�kT��|`�|�.b��)Q��S7�+�����@H�=�5^�1����CoNW��^3��ࡉ^�@�5�����~�<H��<�rhå;=�7���=�7:Xp.>ʵ_[��_C�bV,��kQ���I�4"��wBsE��&��\r+?���4��`��.H2R��Z�D��f9����'�p���5�.���o��J��$H8�S�JA���,�;��3��C[py�@o��עh�I�M>���S�y��U�,��t�;1zl�Yq**RY�@���* �A���$��d9H\B��������&�e�%��m�|,���#$UQ"b1��y�[��5�ppK;���&�\�mĩ�B�ow�W=h�����Գ����~b���t�� �����g�H�-�C��A�<��(/&�z�vf�����w���p��x�f�����'�+^V���?>az-���h�F;�����.�&��1��6�FbhyrC}G$��V:\(铈 w��x��/�0A��u�[23:���'J�A�E�m���0D"0WԨnLV��?5"�nOM)���b�a�M�i(�H��p�.��;�j��?�����e:F l����p$���CR"γ�?��/�g,����4s[v-��3��h�9ǝ�ؼHi�(�~.��o��J�h#�Hюʞ�{�G]o�r���B�RY����G�� '��u`��E��/���h�?&#���1:!�9`��"�}e�w�䇮j���Q�&�P�����|���l�Y�;2� �8�ٱJ�R{���O��J#̕�B���6	�uTX���f�.�����j�3�+���.\���!�a,u�1�J��4�D|�i&[*�� �T��q�H-Z"f��Z9O`�'FeA��AD�|i8v�A��0��^X�]f�����������Ӏ9��@��DY)1(,��[��hg�ł�^4����岬�d�2� ���r��jJA�MQ�NxA���d|d�%��1�$��n�A��U4�A�������R����d�Ы*���	���F�a���{Ý�
\{ǄD��+��	{6�����/�Hnj�t1��o��HF3j/��"��r ��I�2�j�=���be�[ G|�R+� ��3O«'��Hly��_���G�|w|��Z
;��cXD�4#��it/7����o����e$�����o���R0}Y@O�Aoߠ:��l��$���ࠞ�#F`�|�l'p�}#�:�K�>���1\��B�R�����u�%��EzТ��q&�Y
�f��#�Md�|C�]��?�d�+�v)f�`�ӱG�4R�L ��'Ѹ׍��5[Cy��8e�YN5�� ���۔��J��q;�
g�ײ���E�a�r�N��I:���M>�76�\�{eJ�
>?��(K��1��c�������@�����R���5h3�o���LASL���[(L��sn�9�\��t�6�׎^��͡]OW�M�xM�byL�N�I��2��@ʁ�Rwe4`쪟��=/$�Q��L�XP�Vi	����������� ��ۙa����R��L.����T�������O�&���U#�i��^6�u2�Y(yoy�Q�����f�s" Z��`����̅m&e��tZ\n[�#��š�hq8hU�ɽ��V>P5���go����2��M��_g��3Gm0̟[*>U�({�p9�)�H��Wo���_�{�
P�H��(�	m!V�N��� 6�#RI�B�� d#�ڏ�W�K���J���4��-K��-�E�h*���K �ȞJ%�Wg�8�����hT��
F����t	:kng���D6T�������y�}]�����&��Ʃ���U\�y��Q���9L�Sz�k���4�R8G"�����IE�0�V`/o���Vg!j���9���/��T�k��
�}��̻�3̌��3�4�L$���L�>*��"Z����<# J3p=a���ũ<<��3�Jn��4V)�����V]==���X{���΀I��E������<�GL�Mh�/���Hd!0]Y����_�ظ��vh<(���Iaw
N�6�k��C�R>�qn�u�tLަ�WX��_k�=�E�2g�1�ʚ����v��:����0�<�;���PE�H��-���u��k֟Ԗs׵�����G����F�������a�������IX�kG�����8v&I���������w԰��(�'.����'�j#�8�PIAڡ�hR�<��9���u�t��{D�f��R�!J�,�Ē������!�;~�N)$��x�U���Ξ�,�朠�C���^���'/Ȃ.�L�U�����w��g{0��vX�6N{4`��@XX��f����ޜ%��e�Yi�߿R0��v�)��FN��0�ǰx/\�ѥ�|�Z�C��"g.����z=ހ�%A恤Z�'$�`uW�p��5:����H���`kSj����ƈ��o�K�6i�EMx�]�SQ2 /loCJEgǸA��!�/�/h�)�q����k��߅ym0��(��g�z����rvXDB���DRi骯ĕ������ ���m�é+>0��@{Ek<�x$��>�<sEJ7����q���hQ�J��'�g�T��	q�l^ߩU�.W���R�3���[��gaO�xg�7�X̸IyZ�oy�"iq�PV�{{K$�^+���>э{g���.ԉ-��[h�+f������{���{,5�+J�>�C��{1���5��v�Yڐ��8"���!��K��T����� ��� (#���?6�u��_�_���E�,�>r��a��!�8�R����s�RL�}j�,�J�`߹Ĺ�-Ų���*�X��O��3X�����[g	k�_i���
U ���$Ҍߏgx!���Ѱ��n$z���^dJ��I;�������I�3�P�yw]}Q��=n'���F'�m&��rK�@��f���GR�138N~=q{�?_������9��ab����k�:U���0qi�B��Y �u?�y���">� m��8/!�8�����H$O@�u�� ��G�Ysq�@�g�1�h�s��~��L��n�Gb̫5���m�Ā�;v����@}���Qh�H�Ƶ��?���^WI�\*�mj�b�t�r�=-�`�bk ���H'�t:8k�q�F Im5}�d�+�K�_dgZc�Z��A��K�5���F�D���VG��$���u�S�Ѥ�2/��o8=^E\5��=�����U��gNi���[$l��CcY6L���77�M�)ݏ$���|g��q/��D��l�2%w&Y��8��p\�Z�6w��}6b�*xB�؜��u�!�iez�������:1{#���_�
1����m�e���u�x�	�0���]�+>�?�l��kc(<�~v(� ɨ��O"�Ln�"� _ԇgQ${�Q�l��m�L V�u��'M��~�9�����C��ʺ�2���$���Z��Ie��XT[�;4��HzS���J�'�Z�{��x�U����#�I6#�y�=�{��Bi*vج��:qt��r�NK��OHf��qe^d����=xYd��^<�3$�A�.*��Bh�E�����H����_����sq&�mk_��|I�Y�nj�tI/����_��;ʃ�5b ��=�%v���X�l�;4�����=tX�/�o���I�,�#�'w}�����[�W
D� 	B^k�u��[�~�coi�8��n��JT��,��zHs[��ld�H��4��kI\
��p��0����-�AH_������`K����`��� I�4 lӁp��<>l��F;�*�2)������P��F�()ci�e~���T�}�g�!�h������e���0��/x�Р��me�e[��a/8l#y&RB;c���s�`�Ό��t���QyEy�L�H��!2�̛8�����֌(�����٠�ލ�Z���6�>��^�S@�<�u�I�]'L��T::�$AQi��bHr�kܲ�g�ULP�^ԬQ� 3ӏM�~�ކ<��&�V@C��	ޏs7M����!�Щ��-��B`"J_�M$��5��"�K �M�*c�T����Q��䡫lG��JmB�^{$O���-6��-�y`�gR9�8P��Z/!��t6�P���jX#�N��9-=-�m�*�խOץ/�T��zI�\��A�pC��g�����T���fC?x	_5�2����m+"�����p��OK�KQ��l�ĺJ�Jԣ�L�-�/j�Gyr�_nt|��YN� #_"��V� zP� �����Z�bQQ\[%J�"�\~�� �&i�QP$��9��,��;]�ab۬iغE���	s�t#T���:���++�t_Շ����5?k�Ք�C@��Z=���t�
b�=���&XJ�}tmP	�h��~0�O�F�̨͞޻��lR�]��ی���EŰJ�,��հ�C5���{@��V��s͎dJe�ϧ�U�k?
�w�!Qc�H���!�P̕(2Jԛ:U���Pm;�h3�t���B.:� AI�B� �7��3���7zK�+�u��Q�\�$�`F�]!��J]˙�v�IE�(.��y�jg��]��D)����EG��,`~>�j�dwǸ�f2Q���S@e��x�J
�g�{��Rοh��V�3�\{��U�ǥ:~���sU��@m�>�z��)��yS���<6��u�h�n.�FέDom '�R1s�Y��Ca8�Z�i�	��d�'�z
��Ǽ�:���[���Ԕ!å�}Ct.���i-�_���p�	�C<x��%�U��a�0<�b������+�$J���|p�~ �]�6����9�H(2�'�$'���ĕ�(Eh�(�h�]!�����Bv�*��{���N.ةS�]ʨ�9�a2Yڱޖ�	eh�5U�Jo'�Ŕ�NkE������d&����2��^	��ɀ=:ϝ�Ɓ^5LЕ���G��p�� �g[��������T���F�i������Ͷ��D\{��RLƋ�e���{�����C�|�_�����je.o��	�KQ�'�򪴽{�1���xS�6i�D:�`�T�[4�˭��y9��ӷO���������I��f���N�<�Z���'(R�N�Ġ@؟�,���aߘ���#� F�ڭ��������i�j�Bf>��#f`+�h�J������
��*���_�0��?6|Ǒ�"�!��Go��5�d��O���(@GmU2XG�/���[���-�� �?u�ea�nP��
W�{a�BX���;4y)��i���(�������|�*��=
�$���<Ǖ`���s=ֺr0�,��n��Ә��UH�[,��h����(ӣ��%}B�&MΊ���y!��^����M�폚0n����V5\k!�!�R.�-��%j����H�<aϦ��[|�Ϣ�5}�9��2��mR܀��WR�N��?�6�! Բ.$�Po�.������ !I�r:1���sͦ|B�1����j,�[S��H� �^mqG�Ll�G�_@}�s��C0�5��B��_ж��ߛp�[�[�9��M	���HJ�?�4���5� �_��G#S��;Cb����2���Wv2�[L��R��q|h�� ��	T	���H��g�*���̐�'~��H�{w��8�N��$�[���N��F�_��.Y�j�P,���RWD�b��8�K!�g+�)���{M�b:Z�(*�ɝ�ܐ�r���-���~�=3�wd�7��j�~��<v�Dxq�7�h�LG%Cm�����5<�p��s",)d/�s+n�=5_U�
�ʟ9��Q.�g/_��m�|q��C��S���y}cǺ-�Oz>#LS�+�}�孹l<%�(]m����g=qG���H�����X�:��c&z��8��^JU!8�5R��q���@р�,3��m�2 8��+�r�+�z�Z D��镰S͝��C��vJџ�˼|�:�x�h�Di;����eqs�����J��kl���^�7Ծϳ�o�}��j�Ӄ�����H؝Z�l�����Fy����4�f�5��.i��A>�ɵ#��^�����.�<��`ypD�q�(V iX���X�q,�-*^��e}�0h^~��K+p�/����6��*� 󂌯{lB�� 媕�8�G�J��-g��
��" ��Xڤ��G�2	,�
lBV;�Wmb3j4�`n�P
ָ�Z�W�5���fY���^0s/�1��*��l��:y�����̲�.K2����#!̑��f�,%�)�eF\Cj
!�3=1�����X�� �Z�Z~�h~Ot�4�9ޡ����YJd).�������d'}�!�)��z�JQ�; (���1�D�_���ֺLOl��2��6o�k�}���#H������R�sT�dshx[|��7��ڒ��6��f_q�m�D�sU�eS�����N~��֡qE�b0���a��g�L0]����+ʹ;5��2�F@Y�K�~�`�Yc���bm���e�QE��}�5 �K���"�\𠽤��,��ש`�jx�|2B(7�h�d�4!�X��4.y�[u�fU�5T�#���Z&�<�糥��t��Qg�O�{߆�u`W+���`���3�	3���}�nH�Y2I��K}zj���#�v^^��{j$��l�(A�?�_�|�I�4�E�*,��ea��4/�J_�ݐ��Qv"�4�_ʉ�^_�B ��{u�����-�Y�}68��DL!�؍6�0�q�p��g����p�j�n�"���d�ȊvMLq�'��y���x� ����rH���LS��$!�$}Ԫ�S�4?ƩDL}dn�h�ڣ7������t�o�d3���0/ܐ+�i�S�3C�N�б��#��@�'��zR�m����)Tob�lg�9�Ƚ�3Ap��i
��p���}��8ů�$:�\_V����{\4��%�9A�P�$�|W�+�x�\�>A��/]Ck&���@Ef��ެ�ӭo���Y���U�Q���O��{K�qqb�6{[~�!0 T���L5J�Q<�X۫���[��)n=g��C��z���8��(1-�!��c�zF��N�'k��r1Xy��\�'Gf�W���N��B�^N��"���R\��D��LP�����V����1l��K��(j��rT4����}���%���]Z��~X�rU`�T�(����wO���Z�����n}�]�l}��!�G�e�ˊ��W��Vi��L76������k�FT�#6'Vc.�Ã]R�'1���A��BҤ�B����0v�W���F&���N�#��ɦ���]��o�v3�$GԻ5B���x/,\�N�&�2/-�l�M��l@�F�y����r��K���I��i�Z�0�g���~#/��X����i4L݉ֆ8J��L�i��g��ו}X��?��7)�EX�V$)���bJT����;x����#2�[�X�RC���i�El�d ?��j��������IH�8`��c�����}b^��\a��=�]��!�����a����c�g�{�)k 燀X�G�3�:�y��t6�)T��������Y�٥f	�e����f�l_��S�: �x�`�=І����=���u܇��P�~:B���5�v1uC�iN݁��l�g��
�	�e)���� ��sٕ���O���E���)�i}��Q��J��l�d�q�@TGff٥��&��CЍL� R�{t\�{av�W���Y"��Q���g���N~hf������� ��zf�;�4Z���o�<�N����}� 6�j� ���+tg�����a��R�7�DksEg��w&l��%lm�IP��_'`5����-��Ix6X��Die0KB)�+�Z����I���H���]ۆt�=O��G(�x�6$MX�Q���]EU���d��O%���oAj�4����+��9�~h@���!�nD�Q)2�z/���z'�ƪ�񖖅�&�����yx� �~��-1l�J�@�h\���wV��idQ�f�� U@{�G��:V�W"U�{�<�I�0��Ƈf��3��T�O�|���vh�M��D�����hN��A��^�F�|.:<w^n�H����+3�Ô\�r��I�Bo/�D�OCZ�8�d�i�	�)���:��~�Z�w�����k!�b����zU�h8��?�M�������[K.�N���U2�@��o�s�*�qv��9"\�D2���D��O��UV�׺�t#ė2"����S.�SoV��SpY�\��Q�0���"�Zv���ڂ�A&e�ӃY�r����8_�d�":�i��U��z�5��Dgy�4�-Z���}�!��o��
f`0��D�Hi��_}����؀�U��-�pN!��c�Y1
ۯ�2��[=�y�x�IzWp/�RV�|z��;��r�W��@w��۾���{)�Ͽ�4���e<	8�sz�[ڎ8DqO�s�X��k�Kฆ#,�۪�\lTM��������G���F{�ii](�povI�#�0x�L 4��T<�<�Y�qw�>�O��� T�SJ@	o�5�Uj]}_�%�x����&��Wjs�~�+��Bʡ|o&,e�k�X�*���g�chH��s��,/��h�ɇB�@��2A����0=�d�b����:�LDS,��eZ΀ߣጿh��0�F�\-R�R�#�ԟ7q��C�R����a2umܑq<��l����e�O���H�{���Q�^�7�0�TM����E��sN1�ˣ��ϵ�BV��Yƛ0pr�h#s嶉"-a����tUH��Ζ�������)j�����v��HT�a��r@��?��w�f�DE\�6�6F`��[ؔ�_��s%�+�ߊv��bH�-�$���'pK�Sd���i�������ժ��Iq��Q�q�XRQ���~�;�D� t}kx�%>:Hk^�i�w��F �r������%Ge�fx��%�<ds; �ª&���y/n��q�[Cs�t�KH�r�=��)-��՟h9�v��_g��V��v�}�������X�ۖ��J��E���8t�@�i0� 6��Q�9�bi�e��Jmܴ��=gf����q9��quMd-믻�i�c}�K&�.Q��aq��:�]1;GIj_˸��C��u[I[�^�����}z5������N��O�R�&9�Ի�撘��U��nt�(�����)�W�A�����;�ǵΦ�H����R��'Ytq�)��v� FL4q��39G�)z�Ŧġ/�S!׳`MA�3S��h�#�9��J]co��W2J�	R��t��[�����nWN���1و⇄����$?ᴭ��V�
�q[(�:��
��jRp����#CS�&�jP����F�e�xR>�
>�sy�}iw����I��]���7+���K:~@��:u�Q�&��%��6vZ1�J��-sRK�%�c3�V
	 ��q�P�]��- �����!�|u��P3�2P�)v��Ӥ ʵ�6Wq�':��$���\��Q?`�����5��_���j�:|<�gZ�#׼>�B)���ＦD�R���h�ys��<����@آw���7eDd�˶���R��_gƌ��Q��.z�	YN�2
��p�k����k�r�/�3�K3�E~B��ރ�q�����|�� ��Wp���!���\Ki{�1x��Yxߤ��T��)���.�v.4Դ�T��+�]�`���-0���=�������������9(B�ϖ��/���d$�G�+�\�z5>o�
@�B-�dB�h��ǳj�²�桮]5�t�.č�q��	C�@qf��������S.��Jߕu����=n��*�
>4}h�(h��d�FK'�-�~�]o#�ta_&+I����/����pj�Ť�����I*A#�,���<������:�$��m�a�a �s�S\"I�¹�r�L�B�J}�v2���X	�jXcWh3_*8&����Z� -zKb�*�þ��݅�x�Ix�������?�݇3y�J��Kj��3a�dG��Ob�c�n�<3�f�Z��8m;V`�ߢ��l
��\�H����b�� �������"�N�����KG�x)Y]���^�l�7�_<�]
���Ap���� �]l6V�߲m7E~K��F2��p4B|%g'eQ��b��~�\'�
�G�jg '�^Q\QS�6��������G��`��w�o��RG�b��ղY�`���KzbI�p^[%E���T�-7����L3=�C�K�Z�R�L!G=�g��V���{N�Pf��7]Y�֣qxe�'�� �=�eTr���e]���^��sԶ+�m���޶ONӺ��r�2��_�K_k1&<=���w�avюfG�M!�$F�O]�P�v�.����$!o�'��xZ�|5�c�F�~	s~̸U��l���DW'^Ju2wkI�Ɗ6���"�E�`��`f�`���.REXImȘwfwn�O�������8�7s9���'���y�#�>�x���UM�wA]�����_bV���[��mc�	8|�ħ�j,�jp�Դ��_bE��^��@HԬ!�{y�<s;!R�Q�v����M�������^��Y��F�vB� \FP�Ŋ��.EB�.Q)(�4�_�LD�B%�A�o&�bg	䧇j�}U( ̟�E��6PK�}�
jrU:�`BG`��eOA��(UEp�L(Ӝ�@��%=��z6Y���3y]��{Aďw��H6�v�?f�`_�`�Kp��;P�A�Ƥt�4���y�U����k�i��+�Q�4s��}ĐNn���B�g��5i�̺E��p��j�J��B�
J[�7�k�<�>>�;P�Tj��BFAix�Ӽ�<���x������2:2�J�AM��?��5Gэ����Q#
k��֣ ��Qb�P�"���<sA �ru�Ҿ_fK*Dc��6nМl�z��B��7��U�q�>*�oHzL�G��1� c�nb^vP̘���(_���u�l�	�TMx�SQ�3�f Lx��Z�хL]d��k>d_�<i��R�0*��S�ё�c�#�1����f�Q��c\U�L����tq����Ԓ0q�T��Ԟh5vؽ��6�C�w������S����7����M���B��:E"��	��sh�~�5��HO0PU�	�d7Y��[T4����_�?��huy��������O�'��[���������!{�y��<�W/]l��I��e7H��{���E{��+E[1$\��h���v��d��0�I�/b��2�����O�X���_B~A�)��z�/��})zEV:����j{����Ku�$�h��?\W,_�<����3���D��1���|�N��~�J���#W����E���9����9�#,Ei��b�Ȯrkkנ��Np��n��A]hi߾��G�#&�z���4F�Sa���l,� �W�nL0�#T4>$�+ .!D{��N	����|ȁ4�a��?$Pg���a�7# ��}#����]G� ύd�(6�h��)�����Ɋ���Z�������ݚNC�K����	�а��_���,��`��+R=���/� �5s��?�8��tj���	��I�I�7�ZNj��{L��cF�۷���"�%��Hhi>��~����q(o�[^*�.����7�:~~|r]��&�N%���kI�;5#/*670�f�ep������,��C����P.j�z�=u�7#��Sd��y�O,�U����|l�<��`>����q3�`Ϯ��P�O�G��H����;``��DD�Q&��蛤��7h�����A�pع;�p�\�<)�%H���V/�?��$A�Z�G0}D��S~��ϸ\4X�[�'�������oY��F^��w=��%�,BBd��S殱&�~"�ln����\VfZ�>g���;���ۂiWP��%S�hd*-.ړko&�����͟fsI��^DXw�a|����0�� ��,-��|w���G1(�	ԊijL�M���L�b��K��¥����С��NM�V�~�݅���8�&��պ�*Y30=�m(?��E�����l��}W����5KT���z���l\��ڡw[xg�������^���%�mX�Z�>�v�魤���G+R�S������ߴ�3��]�-:�ab�#lJn���˫M�o;AdqE'iO=�ˎl�oOJ����pqܺ��K�u5���?}����:�� n��� �z$L��f��$�\Qޱ����m' �+��s��g�9"����$�;�o	4�����d�,�WG�
k�h��/"�|��+8W[qp@]�!�o���j����n;4����<P֊F�($���`U�t�~d-H�E;s���X�f�qA�i��H�a1�kR�����ٕ_�s*�0�-p��0��h�G��Z�-w=�Ȗ 7�����WY�Ү�9���lн�����t�����V�QAߕ^���luX�Vʹ�=�_�!{��.Ǭ�ۼ`~�Z8�8't���B%N���"ҐSzЍ&݃:K�m�@����$��	�� �7�՛%Q<h��nV���J�_87� �۔�>�&9c���d��Z�������H����bb��|������o"b�qп���.b�
�`�� ��M���˂�ϣ�Ad��J(�s�o<v�~��1y�#v�c�����Ͱq$��프oI�/`�H�+�c���-ɓ�h?��\O(T|(p
n3�X�&ݵ��S��1
W6^ƑL�@�?3䳦��������� I�[*�7���������y-|�]�:���ᘐ�P	GX������6�c���^R/�K�9����
ڔ��.=�D�ޒ� xY�N*��%��+�6W2ׅ��������dWݱ�@�[�jU;�4Rt?���7��i�8И��q!�B~I{]�Tn���x~c:}/�*p �O)��AL�!6� �4
���l9�_G��^3d�L�����7U��<��	�ګl�0�M�θc$��%�Ś�lG�CPk��>�>_����u��UJ����z8��7�d��i�sk+qP^J���uW���j.��ڱ��<E�Ze+8��N?�;��ӟ���\5O�ѣ�j�����W�u#��_���#r~A��mJ���=���̓��Mfv
�fVV Q��󟔂w���3;���/M�E���O�4��O��8����nvH��Pe[��+X�r�J@�iڍ�,.,��7����/�Wc>�̘
8�]��{�?�ܸ�y�k�����qz{90�v> ݏ��B�(&�><)W�^x^w9�%1i�Mu��AT����|l�2xc�.4	��H�M�硧ą�5��|���h�e�j��8��*.sr��샎��@��C9|�*dS��zr�`g؞����Hy������������f���cL����d-��*���>}�`�y��d("��Z=���|X����D�漊Rg�mx�i[�q��'In�J(�:�ȡTl�(]Y<讐��b�#>D7�@���+ �z��5�b���vDX��${6@"p-L1��'1�oi�6�_���G�-��~�ǘZ~��f<ܥ4O�_C����������A��x��� ��	U�=���P���9<BsۊmP�-\[���}�2}����C�i�~�N�L����n�B��G�#�Z��я"�:����y�iM�Q���C��"�BA��N&��E��}�ӹ�Z�ݭ,JS���V��t~�SN³�s�)������?FMB5�}��Yׯ�.�;��'�vQ��nX�B��5��/X�y(*����q���t�P�5W6�����-T���k^:=������0��zJ�obv��x�s�D�E�tAb�����0�H��Zy��=�:V�:��G1��y�	�Q'��_��P4V^n�[����W�2��0����9}��u�-蓞W�Ԓ�Z14�X�i �:,�R����iR)�����^h�*��D'Ġ`Kю�_�� _Фj�`du;0�������j�AG���̤L'PY�!��vC���4lTk���'��sd=�2��'�m�T�	�Џ�|�;���&�RYh�M��;I�e�B��k&о����0NU�lC_@��x���(�<���L�[�����Sf�T�]J�8K�j���r���*��� ߚ����Rt�t�ȴ���o�N�n�?��G���h��Q�5�'e�N)ʧtj�����ȜJ|�iǯ�m'�EW0'ۘ��ʹ�6����1��5��R�\�z"i�%Y0���;X��)����J"7ܔ����M��7%�D�% ��4��Zb�瓩���T�
Eܤ����Y=���
�ٰv쥦k�"y���� 4s����EO�����5�ӗO2J