��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<���I�������w>�sc�˧�� )v�p��}�)e�RRD�\�0NM��Sռͩ�kBP�����K=�xP�K�W�6Y,Z����k��'�?D��;U-�&w����-�lX�A�>ў�zJ'���sHuiX{4K
�|���R6�����

Y�1��խ�$"�A�b4}��߃P�{�O
<�;0��ܗ�\6y�~����t�~� �0�7E�"b�������%�y��̑j��.%Y�b�e�^��X����c0��:��,��8�K�!!�6&���,{���0�� e]�sˮ-\He+#j��ɦ:h!dLy�63����:ڜ#�	�ԹK�U�gzB�+s�܍O�j�g��������#�� �cmMD,{�#�#�T��Q�b�^<��B����v'���Ã�U�7{_�R=Xs0�@o�P޽�������:X��f�)�`���;�Nx�H  �Ou���w���+T#�>��uӦ�
���Eٶ��W�e�Z4�^^��9�N�~5���}�,�h��U��|<���D	@s���G�j�X� � �U�r�zk�'�J�r� � 
��W�.2 nd��=B��G����˯יRg�*�Fa~� �����]�H�u1M)'�;{ %��Y��-~N	�'j��V!���12`?
��>u8g#��J�B�s���u�۳$L��X/]����C��P3�?凙Єm�Ξ�JtB ������^u~Y.
 ՜_�;ի�/���=�U�ͦ5����!
�!��uJ:����3�	�q���l�f8Q��"�<��\{7m��`Cx�`�=��haa<�r&1��'z����1����DX����
[�Y��L��H�7�T�Et?��%	<��A86fuSF�f���OL� =�0��w	8����F�ͤ׺\�f PQ�E0ARE�%�I.Q)4��m5,m.c���W�̝�BX"/U��+�a��|�B�{)��W{e/.�]\��r1�m?_�l6�'���|ܨ*��:�$	