��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<����6��V����ǬT��[Ò��=�Tlu@nA}fq�@�~�U�>��@��mL�<H�p�-Υ�ٖ��$i%M�E���t^��@d�ص3��`�3s�g�%X䌞ǣ�!�q� A��'B&	���v$BKS^1Rv{_�i�湘ި5|�5�E4�x������c@1�#^ߑ�bi3*��SJA�:jc��O0`4��\�0�Y��Cv�p�{��Z[�,u��%��E���.�S�[�*�נ�aTS��-+�ʮ��b�yJe�y�2�E׈tzһB�Y����U3�~���}�F�5~I'Ҁ!��b�]>��D�6��Z��F���Rs�~BP�A�XЀ-d�����F��}��I�Au����,�1�"�y�!2��@ΥF�����8�Y��t6IJ�'��{�S��%Z�����^�h�N׌λU2���*F(�~
|H��u_�j���+����"�k�a���d(�<]ٝ��O��U�񏵑��{I�l��`b_Į�Z��G��0�S�0^%��b���1<�֥:$�٘u�&�hp|d�9y�7_��b@>E�5�{�`�������l8L��A�~ֱl�����I =���g�A��pI/�t����.6�����݋ܫ�TYQf͚���Fm& �9�0���}�t��&�
�P�@[VJ 4�~� Y@͹ݿ�"�/_��?�,���*�\�7�ԇ���^r���o@jK\ӥ#��)d���_G�ˊ�?�7E�t;�c0��-T"��.��xY�(��- ���ۺfقT3ˣՑg��R�.�1��D7*���������(��a�տW��Gj'��9Յ_?�a����}g�Ǟ�Si)d`*�|��ȏy:����ji���{m�����>uV�c��I�� *_�y=��*
�C؏�k�a���R�(>�S�1��,��>b�H�����]����m@C�T�}����4+��ߋ�L)���W����E�F_�J��U���J��ļP��πJ��X᠚v�z�se+E��c�>�Ó��w�^�6��&�V�d�fe��	��A(�g�6�����_9����t���j��v�o�'������sE��f��i�N�y�TY��ί�1�Ee`A�Ϗ��r�a:(�D�?���ԩ90�;�	�,�y':_��_�3��ڠ��lp��W�iY�vJ�c���d�r�A{H�����ܽ���Ds�~���}�~:��3b)�@�����?Ȣ��p?o�ͻ-�K�ۃ^�j���f�??ΰ��ԫ�* 7��R���Ws�������,�){*�^���)nn͗]�unT�rL�+XB7��dG
���G����~a��Y}���L�r��I]j��3#s���kI��_lx���� ��
�	C���};��J�I5t����8�Ó3$\����D�3�6#O��\<��3�D�����Z;�i�s7K@A	VM�#G�J�қ�f�QH�X.�\�X_U�����0x�/(|�
R=�������+��v�bPx�4*CCR�E�Q��e��z��}��-~p� S�X�'Co>Yo��O԰��j���D��.�﹔\����q�"6�O�Zv��WW�_�_l%�:Bf���!k'Ӄss��r�"ֆ��h��1d����EL��]�RW��K�z�B�[D��+��(��U#-�ȣq�\ՏC0S����C�m���#���jO� �ъ�i�z(6S85z����t�lsD��\?�.f�]u:(�ue��E��}���N I�׽�4���-\n頦@��˩�_�:��f���(��p��qh��YIjp�rP2^�W9N�Y$@\�&�]�9!B��in?�J�g�+T�v��!��O	h�z԰r�D��W��
I���Ǧ�Ď]�@��q3ur��:��6��iH�0�<���#\���7�fEI\A������R�`p�`!D/������iP��n{y*e����(|��VݜK�;��t�w�W��
΢h�V=6��+L�H*�Y5�o�V?|�V(nJ�\�/l8ǖq!�b���8�d��呚�>5@6qP���prr��?��}�����Up��"�?\�.b�^@��y�,�	f�Yqӻ�XAU!��D2�V?dP?Cj��緯��;q�Yp/~FI�G	�3�GM���OC���.q�SY��ȶV�� ���I��xE6�S��`v.kPVE
ȅ��� *����H���0������!�1݂%��/
'i����AS�PG����IqL��`Y�(��M.j�5\��Ƒ`y�=̫��F�&��EVD�����s������%plќ��L�8XТ	��% #zں���x�zM1_��ᙄP�2��O�.x}�o������o=��0LU@{E��y���q��~�ؽ7]���C��2.li�^&�A<�V�nM8\��`]���5��Jr��<ZJ3�S���T��
~:3W��J��:���
,GS]��%��7�ȃ�d�7zA����'h|6|�R���~�h�܎OB�o�7կ~�
H\���v8L�:�=��f�Lq��y���������b�ﶮL�v������&<i˿�����!H�~�߃A4e��s�n��N-B�G��f�sx�J�~��Z�~���qU6t-���;>��թ�����bX����@<^�Owd@$�0���}�	+�ɽ�sЅ?� �B[�/5���e,�C�ω��p�: 2��5�j�HG1BS?�i��u���r�>b�yo�/��r��I&'Oe�-U�G;���Nox��r��w�&ҟ>|!%@d�|"C��#�!v��Ng
��8U��cÚ"������ӑI	�9�D�y[Ӕǁ˂�?9�{���*�E��/��z����5�|W��UP�8����@�6�E�g��<�v&�6�
c�[�A�>uE�q�w+C�XwPUf��7ř��0�:�R��R�i��a��7\��A�x������a�2��x�z��F�b�t�ZBu��z>٢�c|_�M7�=�:�ṭ���@�3j9*h� ,enԪOmv�=�+IP�e�'����0��*N�v�Y!K6g��+2����%��[j�������_��9�Ő��]�Y���uh���oyf��v&��-�C�6�4O�����g^���SJ������r�p�5H���#'):�p�����ϥ.�0�1W��p���h�o��)����`��NME�n�5�HH.�UAm�4�SǶ���%����ܘ*�D��"`�����D�U���p	p��r�kZZ�脵'YIA1�<�e��n�<{R*�^n�=,�}������{�|hP�=�Q�(�a��sBʿ?��+�Ȭ�^j���LxX:��&�%�egƢ�x΃h�z���Dx/=57� ]���I`HYwzgB<�!���cv0�?�?wk������T��H+�V8Aq){<dc˂ͳ���.�_�LX�0�Ł�y��"*�zޛ>fWC�1^:xA���J��w�=�/�$�h�����ln�,�Lg���g���{	>�Q@�T��S��G�b;���ڸ�����>�!C�՘Zǹ�rYOd��yuA�e#E�v>�]}{��"I1�@�L�ʥ��0��)0���Dc�c(e/2�ӴI�� )�͕'�U��50nV8'MT��N�ְ����}�<_@���V�z����i3�H�����������6�)���X�������qLr�Ǯ��9�?WCc\�sy���3Q%U4�V�Ў�Q�hx�.������?�uJY�]6d�O��®f�˺v'�$M/@$�a��Cx�9�iT�  �UGi�_}�Sf���bmx�����sEոQ�>QZd�#�*&E"�[�Q�e���Ӡ��w��	�S���{
��I]�l��_F�IO]�U�. �˺��ػ�m��K���t�g8#�}j��,A�t�[��;�T���_����-h�M,�~��m��_%{�JR7�
f:��T����g�B^���o\���$	�J�xh��fo�!O��:|�~�Et�h���/�3��_]x�V3�|C�n!�Ϻ�`L$N���p��(�&��v?�;Dn����ʊB�\��|̀�*%�6~mAqH��q�Vaa����\"M��[)$��S������`1LMHS�� ��5̚Wۍq�/.��ͩ1���췚�s£v������Ԛh��Ӛ��!���|w�`2Kw�V����4��#a�+Eo�n��KS�4�%.��tpQ2�h�R��������R�&g��O���W��3!�-�v��2`)����%��ao
�����<�E�����r���X��;5��q�i�Z;el�H>��
D ���]��@��@��?GMP�l���My���T=y0��q9���_FG��7˾�z�-t�)�I��x���4,���s��� ��䟆M��1��P��g���P�	���N]H���5�Ԛ���f�g��U��(��J{4�I�h_������m�L��Y��;!	�m P��g��U�������"=�Bt��e����2I�]/R�ٶ�$o���K�)8�!��2����;W�/閧|~&/�E�f�M+�I���+DS(��^�T6\fSq���&�� �����A:9zW����2�P���c��j�ǎV,�%�p��X.�y����u:��T�l:��������Ȩ���R���|���Ȧ�S9b�}#~e�(�W��5Бy"Q#�Ѐ�(s��o�����s��l�(HX޿2Q��
�DK}�o-1����}l��"@l���e�È�f�b�>
]V�CP=|쵛Q�B=�0�h������er��c�5a�R�ph�12����b�#�& ���2��#-�>]�W��:a`���}�t���y�~R޲���xe)��2�Q�������XsbN\�M�µsz诨%�eώ��[�"�I5��"��.(�k��-����+s�jp�:NS����7�v~'N.]��OT�a8nX�c��_b�
֓�6�����-䤀_�/�%3MW]b���u+���a[v�D%B�yZ3�M�?����@�C�G	���j�v@J4W��&�� �c2���������%��G�z�B$]�T��Ϗ�}*%�@KϖPx_5��N�̋�u�Vj���9��&jI�Ƀ<�2�X��gF�pu�h�w��c��^�ߜ��h9�a�c�|A�5T��;���jĲ�W�m+�KL��o漏�;��6��^A�C¹V�|F�{�p8z��?��2^2��X��<zL8��~����✽<w?�f�E��$ش��eM�Sge@�Ivf��D5�m�%sʚ�`+j���f�L��_�k��C>�I�VX�{lB5��A�?W��Z<����)���s��jE����ؠt�";wcL�L�Mp��N9��귂�⠹UP��oP�qO�v ��b��ٿ>'�����L�t�Ix�� ����v���o��6Pz�ZM����y�q�6:K�2�Q��0�y��'+4��N��Ek���K60)��I���l���'�زJ�/N_�xv�\��W�'9��w1G�����z�'�]oqk��)dL��{��&(��D���R�z��H���ۄ�vU�tY��sl���8#��V�VʳYgC�#V�D񫪽D��<W~�[[����@�XV�0#�1hɴ*�۰��X� ������w�xf��Ҭ��H�wxl����=�4O�8£�*Z�������!�M�E���b��e�L�<�XD��0E��$6#n�t�wҧ�	._���	�������!�GHK;ЦhM���r����(r������H�fsX�2�ó�c������-{����l;ܥ�L0m�3����Hn�nt��ec��@�tV�� �L�l
�8L��
K�<!M��@!�?���U\=�2�F�&`iZ����2�{���\Bܢ�%���+�f�Z��������dg�KzSxlˆ#$��/���/�:�=	F��]����x���Mt���Qwfa�,@骒�o>��/�#�C����q�U��t���*r�A��������b�;1���O���pД=�1Wi�~(�s`�0�g��|؇��K���f����0D�u�$U�lV�-g�\,�H�'���F#A��7ā�ga���m�SQ@y,M��[1WY$nPdl�G4�l3�Lע�V�i�%���EE�y�+���U�9���Zm�U�t�.�hCh1���9��^!I�F�=����C�Jί�����uㄉ���-'}Bd	=�������=8
�t��?�x�Pr��L?3��0v���D�aY���Yڼ)=�$_yB����b��CR8��Q�K}u��:^�t���Ղ�*�(|��E�lK�(,Zd�ѡ܋8 �p�q��ċz���d���S
�} a��`shJ?��~�rԂ�p�#���(����е�a&9�kS���[6�;�%<��[�vp�,ܑ0����^����M�w��{ËX�D���$oa!�pi�^vDE,�RC�9.~|e6H�d;Be�$�ѝ�5~����qB�Y��Db���ܝ+aB|}JN"��ZFp����9-��Rs�2{�. �W��c�M��m]V�3�~Z�j�u�]�"����\v#X(�đn����Av�)�_�4 z��$ug��3����#T�jwf�Ɲ/�;f�����%�P �Qf�mpm�x�WE#��6���or�v��#	�|�_npkM���P����NU��o�
��~���T�����3e��6��K�-�,�I�>��v�������$ꛜ�2;����M�K���);'�X� :\�ݪp�Q�����tʒR!3�c��uY��S&��+}`�dُ���*c%�E��`� �?I��`5�CD����&���@请�5�FA�E��_������5�C�O���_�^)�+QՁ���q����F��V����T�n��"Ǆ��#��G�s���� ˂4��۫����k�1�z�ݲ���A˛ ,TfaşX]�r���>�0���+.m�v����`�Wg@��U@�Z"�z���K2��L�޸���!m`	5�W9�a	�j���LH�0�W��Ob�vB�K'Yrkmv��Ҧ���g�<�f����(����FZ��������$�w*��;&ҼzG�)� x�"�A�E/`�OG��̙u3%{�����I�~�d"9���Ν��!�췮��D��W�"�.VJ�e�g;$���@�V��-$-\��cwڛ]?S����	!c�u�c>�r8�M&�X���B/�qP
ZCRS���jG��Y`9^���J��cҔ��(��K���o~��s��ӷ[��sm��� ��z���_����]�٫��5�7&kF�{�.�X����+�ha���/m���U=6~�A �����4�yK�&�*C ��j�J �m����j�PHP��v��;���^II�%=�7�z)(i ��=D�N޸��$��z\�@|��s��w�lA$3���_�T�~�fo;"�91I����3�p�a��aф�U�m+y�����7W��-x���x���'�,�t%�����g ��k�+{��]pj���kVV�� ���!e����6�HJ{��hz©�"�8$	-�ƛ�vrC/� WjY��V�g+N�h�:�$|,��Ҁ��	�2EB5B��&������7����I�ǺQ�b�p����4��	λU��c=�a��>�DLpe���P&��p�I� K�e�g3�C�QJ+g�I4��s^my�WMB`$$��_QTW��B�[���L����=�e_�f�0a�n�sQ�S	>�sM���[6�|K��o����
&_P�
�$_��luT��M�Fp��m��~�/�UdYh�dAM���t{����	���r�s��%	6��d�����v�N�g�Q��"�!6I����
�x*��+�����>��ewT�ĹᲸ�I�G��H��X\����5\{E!�ve�j�|> w�3��*�)�]�N{�:��Ս��q����v���ū]�X�b�����bF�6�p�E$,�06�(`�8���p�Ѳ���um�FȲ�h�Wa�@˭S�#�w���^�a i��t�r`K��3�}�o�w�Tݛ���O1�z�ľ"�W��6��i��@��Sa����U���,[y*\c��kI���TN��MWC�35�I&�������X�=��Gc`U9�Y��a����w�m�jJ��^zC_;ތ����{��t����MO;}x�<�N;f~A�Wnp%��ԧ�q.�AA��vy�x!�(���I�"zv������j��f|���<e+�Z����o��NU X�ڲ�I�7g�~ԣ��v
�5�2�;>=�`7E�-�ͺ��Q�&@N�{c͓�h��ޘj��>�jN���)+�Gpb^���v$��ُB�.s��%��7��#f��ƖTW��$�dӵ��Ef�p�,��㔳6Cn���#Z�%��.p|�I*����N�����N̍�� �m���,��V!AAG���ZP�;�}m�q�(�2J>��h}�Q�18j�-�pFҶǐ�]J��x�����3�rx��ZJ��䮗1gq�����];��>O��D�����6B+��
�����aX����h���<L�űc����O1H������Ei�l(�̩S(�c�o��*�I�y.˿�w:5���!��#��Fݍ�rX�)�4o�C���O,� Q#ͨ_�Y���|�j�f4R2)���9�=��+f���X�G~ޚ ��� �����כ�$�t�����H������j���?�Fu�ԉ���(��38�n��̳���p�"���.E)p�4 ��Tng 9�l����������MU�p ��S������Aiv��f���g��������b<�VQ���n�]��uc@���Ui�o�/�	ˋ��=�{/2��P�F8Pi�~�;�>M��������ט��N�Y�ն�4��n��a)BZѫ�Uo¹f�s�[���Uܧ�
�Ү�J��ͺ9�Z�X궮yH놂�� �xT߱"��
�dp�њ�5�;��%k�6���4���0���b؝M)�U�徽d��p��w����#H�A��� 8}a4��Fp.�p���zK�<[��YtS�n�����t��[�<0���W�Ya&e~�S��/�R@(0lT�	��y���mb4��N��M����[�eT8��c��QGV�}��s���i2�ΐBC�\�jQ������ש�M5˜�ۡ.�mǉv��j�h��{�yԝ�a�/�W�0J�w�~�z��%u� �$#ق�D����3���k����(-�%g6�p�����Ѓ�w�4�V�<�)
�y:Do{jńM/7vȤI�2�׹�>A�p��Q�d�;����MJ�}��ܵk�_� T
�Qǂ[�(��{��|l\�q!ե��z��,Y}�A�h3�*��?�n
�4H�6��0CDnG�1
a!oha �37ghR�	�m��E�Rt�u7v��$����F��P�wߙ����/QG�Zl�05�l�*���f^�Ry=8�Q:��[+���.G���:@oE����<�:�*��ٴ�\�?�z��!���.������ ����|E<���@ǡ'LCں�x�|��-*^������e�Œ��2[l��f�=H4�S��h��XN����Z�0P�����Z�����fR���k{��hf{�������6�;x������>�-Ț��gnp��f��-��wl�t�{�~��fo$j�N���+D��� �_�=$�slLT�7��T��B�V�[�Ȕ.>!!F�(��D�E���j>W���U���o�nH�+A#g:���mc7l�	z1�c�V���"���6L ށ"b?�A��;�&]�N�>�>�*z����0�kzŝ
�,0NZ�t�'�;ςf�3��}J�4o��oJ���'���x�ƿW�[��\1�́���H7)�U�kk^���'y���O�d4d6�DP{㜽���G2����"�BB�+�����nQC��h�Vٹ��� CU\MEE�Ofy��2�Wt��4�,��!��+��%}��	����������wS��!�z�hx$�sp<:�8��0DFNi�}Ǿ��
%�b�[h���]���u��6�uA���
�vU���ɚ�Vk���o��\r���|����-�$��ݚ�J��^A�������
����$��� �R�?�d(�32v��S��b�X�E+S����&�_k�y_�?��dÇƒH�jo�M�g_)��P߶3�:i#�1 ��Eℂ�*
����9Bx7G�15�O��{�8O���MEv҅�s���B�w���s�����WRgn��+��ÓZ[iK������{%��L��(ޮ�%���
���Z$��#&hK�qL��ϓR�c7�op�̤��5ͪ�g�`�=*�g"�3�n�S�õO�#�0<_����ɞ�]f��Z���o!�
3�}��YE~��a���f���r��T�<��mA �}--�R�.�4��I۶|�9��'��N����X��_��zx�D11���g_���m�-�Xj�16L��˔�ܩ��ۉD�cBW�Cm��q�1BiO�_ð����T���l��j� �׻��=7��2n�un����,T�֗*��H��{�˞�S����w�#.`�@�k$�4ʯ��-�&��E���d�x��^B6�b�P\[� <�� 
�"�� �4�?���]ϯ�u:Y��]�"Y��b�lÐ���H���_��Q��f���0�"K28��b���d��G�.��l�h����B��0@�r���u�m2��.�&tE`���@�@-�˪��4��e�
`�y�w0����Um�t�{���c�r�Vv�Ih*QP��h����R�����Q2�aA�-W21��2���р�c�b�����q��;�Cl��e�}�tkݾ6�Ҟ������!�ɯ����v�B�N�h�$��'h�cs�U��8�$�8
=��$<��7g/F;���Ќ�Q"�kâW4���o�6���$����M�x2����~$-�@�p�N���Qºr�G�2rWv@��X���ٽL"}��9F�qcY�×�)�*%nQ��ۡ�|��
��(�G�z���P�#��*�5g��aj��=l����s.�$sO;"NC�+�/���A�u!R�%~|��	g��1�$��B���wf�"[#=�K��n��X2�60X��T����N=% 2Yi%��<�~%.R$\x��YPw��3���ʺz0H`��F{R����uS������w5*�\)�3^�_��q��8L(�&c�X3�/���%\ۿ�r��=׺���� ���{��W����-�7��
��k��m#Y 2�L��\�"e!ug�#������*�$W>�d$����uQ�i��~vQA*cu2��t;��jb�S���'���&�oS�u�[�7�s��O����}G)��#�e���V��[���ע�e1�����{R��]�o.�GS�B�~峃��R����+9�+��L�@��U\/L�1��8moe�p������:�ϿV�W����c7�n?*��}��,6�����4ج/w+����f2.�}�n����>��h&�l=2Ê�N�N��%K�
>��-��б6u�P��wi�����v6§�I�q�p�]���Z�&��N5xd�Lz��mT���r5�MW�^����Z��9� B\R�~z1��v��R0:��ؼ�{f#a�aJ�gS]�$ֲۤM����Ә`�J�����Z�#[Yv�����'�ib�!�|�*��i��Rc���9��K�(�N�Z��U�`�G�:4񙭬���Ѭ���z��U�X�dWI�$Ԁi���8)�$C%�`��̧pts��!�W�������K�D�ΰ�o��#l(N@�Ot,�w5�{��~L+ВH'z�y�x&(��4:�eV�l~*���]�:�28q	#��2Ej�"��x�^�UQ�
q���k��Uu����_LyWR��`���nv6zb��`�ᇙ��ȷ���(��i-�l�f���gow&�gT����DǨ�
��7��[����yt �6clA�H�������C]1�.5DK�?�L_LL����IDc>��^�Nc2lvd� %rO¼8���"j��o�a��	���Y��'gֶ_����:-���:̀ɫVw����?����>p��83=�ď���Y2-�&��Lq-����5�Z�����$�~��i�l�Ov�Q�T��	���X�Q��p�:�J1c�&#"7�:��S�9[�[D��ü����ݪ�`��Ymk�����Y�[���"^�?�X��ZUm�n	V�~Hfý���t�7[G ������\�h�!b�r�X�H�L��E�&Ȱ�\^�����{�.^�����^P���Q�=���"cCG�qb�omb u��#�g�r�]�4��M�����F���Ң�QN�L��-�T��ƷC7�-z �R��E����D�&5$�����s��nW4��_����GЉ(�P��}�tUvS�8�K�/�fOQ"��BxbѵS`�NԸ���%��Ԧ#+q`QNl-�XOīi�6���]�1t�,��k���b��#�8����|�wT�_2��oҨ��!�[\���>a0��v��<��)(�Im쪺������ü˖�i�J�A�J��
J���L��ξjW�m��͂�����e��wFu3������9���0,�v�|�����PC#��G�gZ���r�%ri�+z�L�Ml_��1�XUL�j\ff�P[1frZ<"��2�@^F�6�>�_[#�9�=f:�� �r�Բ����
�&+��6�䓠;?a�pr���O�C�93aV��o����9�K���L�(�(�2̦v�鶬˿�>�1�OU�܆d'��9�+�E���m�Þ8�gN���.w�ί\��?_��� ��t���h͹��]2������n��s����)�"e�Nz�k�P�FKv�ҷ�g�=!H���nC"N����r���~.<sEg�������+��4����(_�7kI�8/�5b�0��B�
�8��N��c�ׄ
��}���)�uF@��S�EU���Mm�fS�,�5��
��#�B=�m>�����ws_op����"��ʷ3��υ����#������o��J,�2�hދU���;�乬7�(+.�_\�=�X���_`[�.HϊT���
R�[1�Hw�)�WY�{����R��KnK��.�~�cA�嗶��(��VF�B����e}���Vz���P0���KL	��u�Ep��֌��Y!�q	�g�mP)�}	q� _���S"���Qa��,'���+Ƈ�	p��L%��Vn�}�Y����)��*����@�F��� �G'v�`O���.i��[�=I%����:}_�=�����t�<_������z+��V}zy4�]�]�a�HLnk�w�ҟ��q��V���Y�ÀH�!��]o��c�y�<��6ne��N2B����0K��6�J���.P�E���k�:�$#�J�%tq-�GJb$�3G�]��4��g��ks�ъ`����r�|���_�wnIe3z[~仕ޥ/�Ҙ�,��pG�	�)h4�s�x�vhs6�:�$&��R@�z��ݖ����p��r�X��h�I�ln��c�:�R	�9 j�hm{���RI�E��:9�
7.�N���J�tPt�u�G{Y��o�W�b,,K��ł�CI��[@�BA���q�ߍAA\���#�_���0}��_��4�D^�[����)���.%!=I7h�~Kf'�?b%�W�nό��@�%ӵ�1ɛ%����D�wB퓇���0B@a��@L\��S -��!�
��n\Y�.�6R�ĥ�f��g����	nXu��MpȖ�ż��Hў��񝣎`��g[4��o��v�_L`?0x���?��iuz�B��A��'	.����h�U�R4�I`���eħpgS�ղIg�hxm>V?���^4�ueI�%����yϟѰrA?�t�NC�,���6h%6˒-��Ъ<�4"��%�6��IL`T�f��*I5���&�(9;����t4Yt1�FO2�����������fQvx":(��F�Ȇ�U+�N�2���R������m�~���}+���"�W@��i�E��z'�Cp�%�YR���onH�5��ߖ5B(��X M��/an-L�7��x�i�IJX+z�ˎe5�������`����ȃ�~'����)���,�]�f͇.�n�rdc[>����{�ad��ڐ�����szVw�i��i�����MHd,��30�aDGSA��CU5��)=����L�&�AW:�dO)X}0Bg0L�]S_�Gvj[J� ��
�k�`�}|�_�B%��ĭ�wߏ:Ec�Q1Rmv3�o��I����0ǡ�g��k�c�Z�_$0F@J�!����Xu��>IwB���i�-,�$_�PLg�eH����ꛍ���x�>�2���~ό݋�
0�x��L�d�&�@�z�JIigX�{�ڀWE�/�XnF�;F�bB<�'�6�LE�7����>���JCu<@)��/��n7�e�����:x\��k�E��Y�#R7���]��A��̲Q���s�
�Ճ�m�c������9�Z�R=�-	�-��Z�W�Ԋ����	u�wt�V����ׂ�Yu�'�9�c��CY����?��lEbdXr8���(A�VG{�����^肓��t_
~�($7�hPu�K����p�B3و����e�ݷfl�td!#��Pɨ��5� wXk����}4�H^��z�Z@>�H�>��9���zt~�(��*���)�ҝX@�@I�o��D܍g�Qu cEe4��,�T}�$'���{���y�'#GPe���޼�e1���`�F-~2��t]K?�M����Ǩ,��U�0M�d}�����R"�f��.�q]�;�&�	��G[�D-h�Ӌ�tun��P�O]� l�g=6��_K��7��nd1c�+G��M�w�V
1�Z�$� ���gsQ�̰
����5�<HKV�t84G�[! op1^��]��n�6�<��F�m�g���А2	=�p��vV�Ț�f9 ��lV����U+)��� �]X��iWm�3��f�/t����a�^>��}�pa�{��D0�n���h����]
*��)S�{�i�񃞰%K��q�����J�+F�f#���c��Gl&����#��6���Q�,���H�� �#2y��S�F�_��~����+?|~ע�E���gvG��m���'��4�a�v[�(�DC�� �t�����jGy}II,-�?=�a/?�7?Z�/���	��u�2Q���ٜ�zm5�SYt��9/��:)9����L�om�cͤڗ%�jS��N���(I�S4�&�=z�����9L�<�f���(n��F7���Z���
qC@ZQ���U,�������U��Z���3��;�,�O2���Ks\/H%=Eo�[���z@AI&GSpN����z�@�6�B5��C�-�VDL��!��BW�s�-!B�<O١Ɗ���ĝ_�C�j EW`�n�!.���ciX��o�ұAέ��#t
@>��Q/*��D��Κ`>z|={Ž)�ؿ�9�C�2L򢞨�����VV������]�_�󐜦f#�,��f��}>�ƒ��	� �0.5G���p�*i*^���ۖ�ς]�+���t��P�p<b���+���HW
��?}l��5�������c��N>P�G�P�����a0-�v�A�N��:�*cs$�׼B��fwu���U��cC��#%�'r�pi3D|� ��R!� f"?f��Z�"�+fs}I?]S&`A�T]��p,��@���=lV�,�e�3Ŏ�'�&�Us{!�V��X�'�2�ԟ�Y�c���=�
�^vؠ	:��Y�m"2�K��s�PM�����ݹn!��ӑ�	�1u���]�ʭN�ȹPP��/�*/�ʕ9����9�C��TKF�J8������A�-l����C�D#8P�)�Ŗf�f��l��іAyP���i�E��o>e��w{qY�~3q�����qF�n���4����嚐��4��@��웂�HKQ.�c�8��!l���V�E��^CK$��	�]����7D�Ա�6��7(҄���#0�T7����Uh�ս�_�gĺ�DԤ��������ɾF��8Aɼ��jЅ�U��_ȁ��eتp�U����z�ǩ�/S� ���7Pa�Us�8��e4�P4r���p^�r��L$�>q��{]n)�W��O�M��WY��ɂn��X�ҥW��z�]�&:;3�ӡ.mO�b��;�3�=��m^�B�O~G3{�J�"u|�>I~���\6�;���Y�3��P����^�F����^(]���m}�#�8�c��|ڊ�M 1�u1�_�|��!o�g���j4���鋷�{�d�I� R
M�a+G��A^�Y�>)! �B��ԫ�^�sǊ_�:���a,�Ó@}֙s��Yh��k�-��9�ק���̮�Mq��fV��X8I[���w���2��v+)�i�J���8��i���0�Yd��-98�;z��AG�i��`	�P�j ���Z���H�l4El6���&�p�Eby�D�O�X��G
e)�� NNr+� �59w��tj[�V]�?������i��W�zV���n,W���%>h>���@����}��i/�-���aCԖ����U�Cջ}˓y/+�W�Sl�G������93b=r8�˼".����$A��!�"��,��l��v~+/�k�6�0�
u���'-"���~��t�L�cI�a����(~��U�^(�y���']���?Z��~a_��D`1�g�� 2�L�d�,8�������&�i4S�&/�d�G��� 9BV&V���i����?.hR��!8�i����`O��Ԁ d<@$Wis�OK�U*���!0K��rq�Z\ۊ�΂�w:�4��3�#ơ,��� G���ۼKbB�<��A<!���1`A�%K^�/V=D��a:�p^�8���V�J!)7H�XIs4C�Ġn
���b��$�̏Y�L��>�J�u�}�Q]��'m���-F��'�B��������σ�S��TfGшp�u�!+@&�<�I��,����&ųK*3�x2���A����X�t%�0�S8��B�~w	�~*�`��Ϳ��V�,<bJ
���	ʄ62Z���r[믅㔮-�W��c�������E{ǜ�&��uz|Uan�����Ra��ro#?��Td���)�[t�^6%��tW4=m������h����1����4DЍ}�ץ��d"����A��!e�5�w�1���Y��+���uj���(��ͅ	$z+7�t.p7�
�I�K؆�C�IPdo~��"��אـB�l��y�F[6��!�6� ���/Юtc�.���%�=/S�ݢ|���p�|�ڄ*�HS����v[�@�O�W��QcF0�K�z��dT���a�
���3"Dx������#�D/�;,
�b��Ы���.�2 p���>�M��U�0��ߔ��1���טs� f+�i�o�e�.Y����A���ku�jo�4!��Ə���!��eVN^�'���NC��E%�q���A����$T�H�k�N���ֹv�S�_`H��1��s��xڵ5������H�����9ce��쮔NY~-�IC=��2������L�#�{��&�?�PY�l)�8"����à�P(�&h�F3 ��P������^4#d4X���ēV����9��3a�K�����ϕ�q�Z|��O��s� ȭL��������9+�>�;	��c��%U��r�]h�:�Q,-�|!^��o�ҽ[�/W�_�n��&��S8d�@��<83~�V �EK��r���%B�W(�I_�;_���{���sL���7���E���rCm���7.g�PgYQe�.�S|R�曖'z�0e���,��sձ9��Z�������V&YO
�����R���93����$"�O2M�)Ca� ���a��P�Ycz\�b�.s��F���m ��
K��u�|��.��I� �KI����ۛ
���B6^�q��L�aC�� �g�g֬	7B�8����zs�FI.��SĲ��̠p�[I#G��Z�؀��I�mT�*�
0�{���s��`��q?�����T��T�����f��4>�ӳ�M�����S4 �0b)�҉�?��P�?���J���d��e1�㖄�\
���2h:�,x�pc�dM8\JG����ޏ���δ}���I��G�f�����Y4�X�t�A��>����Z[�:uj�R��1�37��G[���Y�"�{��I��n�2JF�58n��N:�go�X��҇�	�lS�d�4��#E�k��QA��2�E'rA�"4aD,'7���Ԣ3�i�&s�P�B��4�@zQXr�L�'��ʀi����a�z�p!M�]N���*d9��L9���:������){�;o��Ǟ"��C� �'�I�[�6�g*�d���M��@���uųC&Q�۞�D��/��z֘jl��T]���]��sn��H#��9{�Ђ>���Ũm8�s�Q���`D�K�:��uؘ�J5r4o�#�c�n����	���S�e��G��6w&���-p�0[.*���	LI)��l}��j���vAeB
���+�KWZ3)F��Z"8�i���!Ir=.i
:asOãf	�ߥi�6�۹��_���
ƲZ7��)��z|h��
Y��HyX����J��s�fv�g�;7����4���sf��y�D��Lm;t�X�='<fH~�<qv��\��-��o���ıѸ���r@:�cj^WO����vh&�e:6@�%�ToԜ���=-O��xX�Z�5SY¹Pd����qo\,9_�1P԰6�_�$�HBv���x� ��r�F�|������Y�`F`��8?�v�e�M5�{08�nV���0��lY]Y�K��in�w��i���n���K�ܭM�F[��[�T	Yj7����N��7|R�����j(�#{��pU�/	�<>���8ුI3�7�6�)N4WՈ��4�B�7Cn�#Vb��;^��h9{���Ulp�izuEDW-?�凗!�OȢ�'��wO?�(�Z�RRfL%�W4��G
B��E}��T�?2z�4�`R��
�Ⳮ���}]>׳k��?[ޮ�L��G`�:�[)�*X�%c�0x�o%H$����NB$O!r���{?l�Q�&A�;�4�o] 	Q_bd!�W}��ES��3b�iL5�[j8���:?��Ǉ���o�f��n��ϱ(OQ�������s7H��0L��I�O͏�h��}�x��~+�c��ǭv9��jEgi ��j6��(��Yd��t0P^���[�=g�Wr�1A�>��.WSk���p�h,�O
���e�ਕH�	��.�
U����@R���u78UЌ@2�GdN��/u8�G�������%8r�٦ �
�G:{vꉶ>_�y�����U�ꚺTz���2f]K���z�\��;#F/_y���Z
�/%V����b׌�����Uߗu΀^������~H4����mA�s�Em���h��'8G�^��z�u�*�{�rh�;Xw����.�!�{��n�Ӻu#�<X+%��ou��p[q��.�os�@�a�a����pn��H`�����Xw;p�*���5S������\�R,zI"����O���y��DN跔Y߆�h�Ր]��h�rCh�;��[�ѕ	��k�5$�:�Y	sPt(X׸_��o}� >/���¬�+��)>���n��$��TVT��14u�8��4��'���ON���%˓���G_a~"]�����6����@c��<��e�M�N���d橥�5?u\+�H��Ƭ�~�E4�����D^�D!d��߮�� 4�D�Fub��Ƌ/��HT��5ӵ�#U�U���X���:�[k_�В����@�Ead`�8��u�u�����E�w�O�Z�k�<�J��{�$�Z4�K���7�y$	wTf����	N��K˵+ө0C�+��	�q}W���79�����]f9�~�|��q2\n��q�l߳oЩR��z�L��?�?�̆�}٩ƚ݆:���\
T��"�
v!�v�/��	�+:����^�+s94#me�:!W�D����l�.AH��Y|����*j0�Wv�k(��jP^�߰İּO�&� ��ᆌ���3*�'���D�Ț~L"-�e.r���е.|�L�mM����{K�=5G�V��D��Ip��}RcF9��ݥ�[{i)@�[M^��9+��H�Z���J�B���'��7[,S��d.�Ê�7�d*��/�"��痳� %>j���5P׏UR�D|N>�H�?�:G_U�-Zyj6�Y�+bMӁ����
B��&%�1�)���Q �ƷA�u��eڦ�O��Ϲ�1d�6�Y>F�AC���U�:e���Έ�gW���o4gH:(�QʮC�.�#�Q�h���b��l1�Ja�K���
4K�̳&�aZ��o�����h9�?P)bG��j0M�����&Ƌ� P�,��HZ����#ֻeq����C�x�>��H��[�pۡ��f�N�,���	LK�	#5��aa`��)X�a��H!�r7[Dnղ�/h�������AI&W�/�zNe�סg�uA����g��Žv� �v�:dv��z�n�M��e64px�q�2�~U<d�� �H9�L�dU ��m�v���fg�Jy"�@H�jo ������?|��gU)U�`פ��L5��&���&��:	k��-,��<X���ݲj喑��.w`��*,��ȹ�����*��[i��3����Caz�Ѱ:X�Vܺ-����L�Ӌ�v���N��V����24{�'�U<bb�^l#����s9���sJ�I�ArŅ���]3�`��>�ltT�ڋ�}�s�T{��gS��nce���r�3�Ap�
��`�]wSfݵζ� C!��ǌ�.C��NP�G��=%w��箈���\��V"7d�e(�������
�w

���&c39�ꂆS�.��O�M��3��'�g�/c����K�&�-z]U��2c�?���a�i���S˵E��Zԋ�:����xc*&""~z�Շc94�o��c~��������*(r�Y[�B�d��T��2�-���Tǜ��/�)f�)Z�\�F9at�H�(�F5Q�91���
zT�_�^[yK�\�#�`_J�qX��	��N���e>f��G`s�f򇗔B'���mE���jq��6�ӵ/�}٦�D�#�y�)�Cx���2�!�Ծ��*��,rud������ڠ5�"ݪ�T����X^l�2�۬�-k���Z��=Ә�3���%h����t-����8�R�S���e���U��D4�xz2�����Z.N�
)w�z�q���iG}@-@a����)��ZI�E��E��R�.�6킀R�5�ZFE)h�d-U^���UbM`?A�O�Mw��X��g��M-�l@�'R�d��Cz1�rJ�+"�yP�]u:"��T��W�+r�����N"��0��"WР�aX���������R�̗U����J.��:ݖ�ȑ�u�4S1�8���>��W6]믮���Oy`���jc{�K�v���٪�GW�s6�y^bc@ ���漚�!��-u}��t��q��b�a�jhS��f~�h�������]Ƴ-h�	��Q���B=�4&|	u�,lp#0��N�'j�������=i��$����Kf���L�W�KA��3�ۤ_��&qg�&�x��z�6N��/����p��o�;�G�Cb��g|��E�x������="A����/�^u�6\1.�+�(�B����d}o3j �YP���'�\v�b;n2`�8i򙺒���D�U`��/�e�F�C���N�n?�����(�y�Kd'x�0z<�ÿ��|�.��]ƙ�K��Q�|����T�i�j=>�jA�*��(��<y��+C2o��r��A����Q4-��ٵ��E,R��އky�I�x�eE���C�9x�v�{��贃��кG� f��G�h�ݺ�~m�l��?��[��<P�K<$��bI{�s�|��&5�f20�6���Ÿ̈́����B�\��۾=P���������V��!`f�
��jK��!��&��ٌM�6��|I�h�����d7;BTY�������N�ş�����j��]\�b��IY�֍T���I�G{Zƨ����do]m�g?���]�`��<�G%N��@U���alqP�n����$�ecřj��!��@+��9��Wkƅ�~�Ͱ�t+��z����'x�X�-K�u��}3�lPi��.Ik"�O�fø3��A�F��y�l�)%�75���T�O�7�����P�&�-�TTH.*�=�yN#�{X�i����r�H߽� �Q�}�"��k�����8�Tb��#��*i������sU����p5{��y��k����κ��Do���;��w]p �|����ߐ�(��O`,5�4��h�ǿzK��Y�OE��y(L^n�cm�R� X�a���!{���p'��;e)Vlt�"��^�ЈO��M5�h�\JŰ��s�����6+i
�5��@C
����?z7&�� ͙D�"����_�}Y7�.vg�z���s�U�<��񧾮Z�:�<m=�w�P��K����m�U�.�f�ԕAL��O��,g���2�u��X3��7��r���$��P��n�1�>|�5H�[��pL�H[��g�M���-��*̶�7{��p/R��p:��I�o����`7b�.�d�)�z�����g�} ���vEw�$�/�G{\�Sg�v��u��|%�gJ��}���F�$�7A}�=#��Y,t�0(� �g8�<��o���?-߅J�<�6m]�êmr-�P� q�h�;�[�$���h�C{ο�K���E�H�d{=S���/; ?C�9���(��
 S��QND�Q�F���D��z/�O�#��O���`�����/b�'��#m�X�혒KG����w�U�|2 *���Fu�tEްς>�>=iPo��u��Z���"�W��G�B@He=+[{��D��+@�������l�[�L��V��7�gn�6��i��8��"
�\�,)���<&��nM�N�ή���V�O�#�7�ļ�胧7�Dkg��H+A�rӝ����MĘQ��lP��<E
Ԝ���%,��j=]�8�Jr�YI�7?捤?�0�R՟�-���o�へ��4�H )#��쵾/�V��6\�¸��թ�*��7"%U�2�Вyu���/��X�S�w�W�^��q��84�_��ZXl�G�*t��f4%_`�=h+D��+����s
),���n ���N�4�&�(�H�{�cf^�$q��J�K�-����Oc�%��F��T"�Y�+?۔�y�(~��\�V�������W\�2�'G_p�E`_�������qѣ��SJ�(��Eۼ�ٚC���Ʒ+��?��0Ab�S�������$'i�ݧ�e����?��PeA�׶����[��@���[���2�J�+9�oȅ/�#�E�����2����ԏf��<���\�G�����s�8�tOa��%uz�ܒ�W��c�%l�W5���+	����d�#��C��~���+'����p���6�f;��dv���l�!���b�9�5�]�*}����g'uq��<��H�zF-X4X�&��ʃ��Cv�;⬨�TI��')�2d�4����W����,n�:��� ]�2����7�����5n���h�)��F$9Ǚ���� )�:Ja��E��z mIt\��`Z0W�<Yn�p`�BSy���nc&OB�xt���<���w�HC�C�E\�����BDQ7bv�������p��24Z�x��7�|H��Lp�Տ���Q��~/���W�
�����W�=���c�n�DY�Pۼ3�
���j=�驪Lh��w����>��"_��j������/�Y�k�l5G�)L�o��-TI[��G�ͩ�s9ʠ��2�քg����X��P���*�>�R`M��Al�u���;%7��7�������.�Rm��a���e���y�*w�s�E�UI�;�Q��s"?�*M-�l�/�����Խ�w��1W��lg��xr�4���ICM�5�+���Q����bԕ�M��g�̈́��%H �d_w��h��.�#D���@�*��'�g1���:j;�12��I�%�ȟK�mQ�)���4�]ǟ�9��9�#�7t�O&�e�Z�⁨�鏈f�����A��,<������+���@���+�IKu4�Ҫ�#�@t���J���ɺT$v�9o�g+��#���C���*�ݟv<��zO�5}y7bK;L¢,�w����b5h��p�|�^��z�=*Up�����y���_S���ȗ�{5�G}
�n�4P���-5�`6�Wf�����0ɰ�F��Ӄؑ��GKؙ(Y���0��k��1)�4��	���?L��M[�t��)�6�(���GZe��4���N]M�������Xfb,xM�0o����Zt͝�S9H��U���ŰЗ�yhߐ�;[�r����Ha�<��=]��

�T���ڀę����+ߞCσ��~�u=��'Cq�oE��w��>]zZ���V�-~e'�b�!'�q��F/&O"��*���1҅-s�;]�t��i#<�gP�LDE�^�����m�9���R�E�c��V�v6B�3�E��g���4�4jyY%����jz0'zz�|�ܒ��(2�j�����^�g.��q���՗���'B0�[� ^fx84�#�7v����j�蓩l���z`�2z)�pHm-���KP��1�ܶ �dE:Xr6HX�o�����Z�I�Z9�/�ݟA�̤T$��e�K�d�����"＆qmį*|�S؜�R�/4׈��S
-�5CB�xg�$<_���k�����
�pZ6�1�z��B�>���� �ζ(�wI�=�Pq�1mǭ<ia�ZW��F)�$��␢�6���V����
��0�&�Z{�\s��Kie��:���l�>f�ϸ�x�w�ݻW�۩�d�Pn�J���BR^�mW��q93X�%t-��}���Q��$��r!A҄�|�Qf�jS?��ӟ�u1������S5���A�}MU��Y䓐����"%�m֧<!v���gm_�Ï> �؅�l��#��X�c�>~��K/�v(|��1T���5��@�Y�Ɔ�M"�.���/G[�Ly;���m�/7�,m�1d�ʅ�u�����-�;���m�@�L��1L!�Ɨ��WB�A�?��j�� Wua]Ԕn�:���a'$�u'�ɯ[�{�55d�����?��%�~E�I�":,����
�;��\���eK
�(�M���`X�-�(�ZU��Z�N�ߊ=�Y)�d�K�'��u쭚ث�D&y+�ڗ2�%"�C�^(Ü�HY˱v�e���X�!�U�u%��0B�"�B�4KB*OJ[7*ưҌ}Vڻ�O,I�pID�e�獊�-�0N�Hc�*�'���Ц���2/�
�_�/�P�x�:��Ӹ����K�`�km�Z����-����R����J>�r��b��4ȷ�1��/����J�G��"��d虝3Bqgn�,.K�Bc��oU9��.�_=�#����dӟF��L`�
*�L �nw�$cl)��Xw�l�EH��^0^�n晐:��B}_�4eԽї����|��*�LM�j����O���xvt��Eǌ����	�GO=(ZQ�!\���]��XQ�8��R�ccwSI�*n%���Gf��Ǝ�4� HBр)MOl����d�8�#'I�M0*E����!������4���R��k���ߩ��h�Ύ��9���Y�U�
Y���]G!�ڧ2��$T��1��OCr^����ϰ.b��|2n���C�j�ml�g-��Ǚ�A� ����ra��WI�ՙ0�mW�Ӑ�"N�p.7z���z�)�)��P����B���ˋ~ⷎ�-c�P{V��YSk�̕�u�K7h���-//�y����}���`,���8%����CS�¾�k`w(��`l���	JDɄ�fz��@c��}�Kr����a��S3o��_�ȻZ��PS�96��t�����xr2������K�!����]�V�^�/��?X����&�ů�`ҠV՜����﫩X��3,��䤱�	�s���xㆂ�����1��Ֆ�r}r٢�<2�e|�7UcrC�T����K��y%4O��C�0^�Q��.gad0��54rv]/e��aS�yet0X#�6�Qԕ����e�K[��M��~��Z���Foݡ\�y�2R��s��G:L<�V��pNG`�/`	�R�������f�w����n;�H�V�a0����v2]?��4�1��(�Is1���:H�`�,���=	'��BMY�\С���u�4�֩Q�x�Ƕ�vl���dg����d���Y8݇h���Z8�a��[�bUO'X�>.�EB��n2�1L)�h�C��4����_ޕ�v��_�gH�-����y�&���K��x�[(F��$fٝ'{�`TR��>��PM�����@Ce�����x�ǟ M�ڤ#�9�S���)l
1���OyGN�����5��>m�����qh���	)�!fZ�LVeJ��Z/�dP+�1e��t�S��R$%k��(�@�.,������a�ſ EH��[j1l�ngm��`���ӳ�uH���@��,����a<�K*],����Q��-3IN��-��W�d.�E��_F����9%�M@c�K�%�k�Yq���A�Yt��S-d���(��x���h���.)f�t�˂ m[�i��?�˲�-%�Iq�]�hwC�S�ɹT�3,�^��Tx�L���ӹ&�N�)z�6Ϩ͂��������f�l��#�1_��O�!,-ҕ�'.,���[�������ۍԫ-Y����z1�!��?}XR�a�4��!��,Wi�ͧC�b����d��������=&�x#9�0f���[9���4yG�����g��\���jɨF��f����>.�tτ<���	s��3����9vj���9haU6F��m� �w��2_©n���8�Z���aB�W�� �f�%���^�?>�P -�8 �)3�3�'�p<s��(,꟯[C����0o��6���8�)U�C�% �QzhF�mo0
U@�+�0*��3�.�v�k�'�Cy�q�E9�8{|I/���YKӴy�z޾ns��q��x�I0��Ѯ^�^8�5��{���@hw�;���D��<�ED6��~������0�NcE��}�`���3�&�OM�ݨ� FȮ��$).��x̉��1�6(�_=�A_Y��]n�uv�	0��TGX�:"�o5��gM���Ò��vF���B7�[U��xU���p��C��\̚�K�/�6��v갇�j���O�H��Q��~�^3�Q����1'�
�ڍ��<sC�,���Ȓ��Ƒ�L��v����'l{�jt1؁k��u��Z	��?��Hж|�iaۊZ5c
^k�d�pW�� ���u�r��7F׆Q���hH�yΙ���U�la(������Hq\�hC�K�{��u���Kf_�ѡ�n�k��'Ei��_�-��]�k[�2x��G��Hwׄ�L����^��ی¿�Ӄ�u>١H��9����'񞐓�&�����擿2p)�o
���R�5����lֶ˓�one��rc�oǼ�Xo�����,�ua��n���ޟ8R�f7S����оX�or	}��8 �o�i��#^�P����JҒ�'g>T�5�R� sB����,�Svh���"A��,���0���A�y�����19Ѧ/b����'��~��V����D�71J�:�ȱEͫ<�eC}�G����3.��_E��2��*�(Q�يrH��O �����*䲐U���^e��ʢ
�b[�^P+��l:��̍�����Q4w��RU��d����8I�MNR|p���T~�d�z�8�ؾ���0rh��ܻ����{�2�#V�����}9���@ae���ODߠ,��z9�r��8�P��8b��S���HN���'��C���%�|ǟ�X���q�k�٢لC��8�9Nk��T�wJ�O����Ta5������ �CF�ڗV�}Ԋ�f��E+>>tz&��J��h$ǆl�|..[�M�B�]{b�>c�=^Xً�[)����T���c�O�r�5��Xgo���l�J��RG�H?"�^�?.���!o���vq#����ⁱ,=�2x��Z��D��fּͩ��l<�p[P7'P��\<�-E�"!	��ѧ��1�.c*.��[lY���xy�ܦVkt��<ݧ2�q��:r�	�����Fɩ& ��&��y�t�֑��q�4���4��M�[��c�>�=�y��nPZ��!�S��ّ��<�&l�-�*�H�W�@���}4�+�v8'�sYx�����o���dT@����5y��-F:?+�=݉(�T(?��i�H�Q匓��ɞ�)��b�p��)���8�7�|���G��q��@M�b�hܪ�)����N鸧�m+9�I��W�������u&_@�.T:���3$�3+)��̤f�]�>�Q"g\�Hc��n$�D�5�|����"������6������Gvp�e�cԙKE�� #e�l��s�3UU�-�$���)���{��d��VC�����.g�N{��itqg�؀�v�'��&)!���p���՞�0]zU�@����3&�B�@}[�"��	�&<�w��C$_]��;��J�����|��u��ű�m�I��J�kG�0����NM~����o&̷ţ�v��S�	���8��)K�l�%T�N��Mؐ�T�{���*tK$��	g�І�;�b�٩H X`
�K͜�|_�zV��.�o��ѵ^�Ƭ�&�3�m��q(��ܰ]�/�Ej�^�k>[�ҧ��IIB�ޟ�ǝ2�&սԤ�єx����|��6\Q�Sڗ��bi�Еx0Zì��¸&��n	a�}k�R�-`t�z�ߥu/�Z���먓