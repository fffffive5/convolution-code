��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N�'��9ۃs�)n�bpJ��B���`�h�v��>�R�D��ɳs����@EvR����s,���?�)�|��l��[��-��i$��ז�����y��(L0.��'�9Xq��ۃ�G�\zK�r�{�23t�p�t	F���uZ����Hؑ���8�9��6ᔜ�@�!�
�w�Q�뙂������zۘg�\�R5�᩶���2$�@�@n�b��hT#%�!iGl�w��/�s�+��l���@�(��{"�F�ٌH��/��QC�so�O��F<R��g������b�V��;��+�v�7<�%�X;��|�j�Ŵ��?�ȸ����9���}��� �7ڄ�2�DZ�� b���Th��ޟτ�FH�%zG���T<fu�G�+���>5�2��.��;Tgϴ�@t�fD�9�ަ�#!,6=��\YW�������>B�Y�]�:kV<�s�W.�ك	�^��:���G�]5඲��>������ݗ���ٴ�A+}=�<*fa�?�|e����i���������76]*��ǹZ�m�yf���K��Y2�%�����mLP���4e~�w�uv2$�^R���}�<N��~P^�S�.T��B����C�U�b�{�JÎyJ��*_�b0p�M�����r]&z6��BI��#bT"��cvtx��ʝ��EI.m*��Ֆc�V�{jd�L`^햼�*ѯFx&"Ⱦ�;�Q�u�]�LT��޼���tw\�S�>pq��$.�G1m�j�0�A?C�d�5`�����4�
��R5���4<c����t%G�&ʧ�܁�4���9�嶶�`t\���ѩ��Ik���R�%��]d�S�m�O��j�$�f����
��'��nD�Ԥ�6xܻB�s<{��O�?����5�C�	��𦼸g�k)&9`�v����l��=��2x��
��4PWa��[=Z\�e��*m�����4߸ZYϻ�P˜9b�NtS u�c�/�Z�h�^�eQ�>b
������J{�'�j<@�*Y�H�\GW�Qy﬜@�b�o Z���b����MB�X�e��b���s� &�8��E=0C`���B7:�
ԛ��2�I[Pշ���I�R�  U8�&��yb?O/��{��G����oc����_u�.��F��T�lV���I��] ���X5�>8��X�k�ioo��gUKK\E�zOݨKPv
퍧�^�K~��B{�����u��a~�H�R4�]��Q	Pr�R��E�q5�"��3!q^���
�O���N9�0�����Gh+i;���֐�7���'�|�ؔ�L�:���J�i�I�ϰ5�m$�#]gO���r ��r���m\�������@�^*��oڎ��e Mx$*@6�a9��
=����.;�N(.��oKS��v~u���T�x��z}�iINJn�ƐW���*�yG=�9�z�ǃd�]�+�tX�"nBuK�	�,sĊ�f�zuq��Gj�{��$�]��IB�z�a�L������$����dS�i)x/���{�D��
�C�l�)*����呚D�5� ��7$|�&R�������/�X��<7?_��B|�q��Д;K��;D����%��#D���Ѿ.-kvR@��	�O>�I-�׳a�=2�c��_�j����\/l��q���u@tFA�W-����Z_*�m@�������|q��M �hH��SO��1�QQqr�t��s��q��		[e �r1˾[��o84�
x�XɈ�b�5~�.9���I7fw�.��Y�3LC}�>��k��`����([i-E	ж����`�,��Gة\��Ζ5����%R�O8US�r�H�Q��5Ŋ�f��X����r�[1��mr�L�������>-��5�=$ibA�_ZR���ɳ�	�s��ֱAg|�b��!�E���]����&|�nJ�
�|Ei!�-T�x1�b6��V�V���:�T"8*��V�/7�=���۩ ��ь�ܢ�,���o�<8h��O�tU&��o\ر�X�^�Mxv�SnQ�\����I$I�6�2���E�M��y��E��pK�>t?���x��������k�e� �U��].0��к`���0����J�l�wҶЄ��g��_���ܶM���+?w#���_5����t��Q�����k| f���@��J���GZ��d����_��\�6u�۩!N���j�o{���8_JE倎.{s2������eX鶱}�ϰޖQ2�6��G�H�+��u0�s����*��t��^�Q�h}c�Y'i��/e��$�|j3[��Z���4����@Qr/rH�����Ksw4Q��,k���T��qH!���W���Z��i�E4�RK������:�����[�|ȉ�I����t��T�\˩�����w�O#FL;�={���5S1�0U��hF�+�V��^��,�_�KB��[)�3�H�O眊ќR�Z%r��6;;[����i�P*���b�E��2ѹ����t`̍�5R!aK�]K�.�l������^2,��<Do �>�l��ة��aa��h���[QԿ�0�9m���`�L�F���e�N��e�&��CD�)�(j(V���!S3
��x�Z����3A��dl,�E��z�(�مڹt����kt�s���\\��r� 
�I�%r@��6	�-��7�b��M���G�������)�Ó�)w�IS9sKAo���$�i�ZAz��i�����̨��S��`؁����X.��G�5�'r�
���S��,$$+%SğSH��N�2�i��?\UXir��ݚ �u}ɛ��&�����&���!:B���k!iZ՝��`�V��������;'IfET	�T]+�4�c��32��b��y�Cb����+�Z��U��d=H����}��k��FeFLGݼh (e�e�uU�����h,)��d`0`��RXa��_��� ���vd6�h\_�N��V2�@�fI��,=\Y �K�Խ����61.�>3��C���kp����X��!?/�����e1����F���6� �W,���;��8�h���ZL->�Yp�6h���V�=pp^^�\�3w�� �|C��&�E�H��U���AR�6�M>�۬I��	X!҅�$GŃ�=-Q������r�O8��6
5{���Ś�%[s�M���1��^�ol��>�c��5�O���&8��~��+���zγ�e����&Io�������&b�I����^f���4��:����{4;S�V��}M"��؜q�ȩES�C��,K�Lɮ	��y
o�X��tGผ^=j�^(��.t��_8�=��ёN��!g�)^�n$�F�:��L�IU��N���礓�#�Q�aq��~:?y�B��"O�p7Hhr�nW����ґ�n�D�a 	-J�@��z�;�Ǎ�s�hV�q���ڳ����hS���������������=dƟF��4�l���1��B����>uG�<�����a�T#m��B[9=M��q��g�K�,��w�=5ev*��p�
y+�`�>���L�95�EQ
��2ajo�Ƚ��t��-X�L6�9����&��w�/�:�~Η^�A�������p�=�#+J@�ᕲ��쀝���z�n�S��8L�=�0o��1�U�3��&`��o�aw��u���X����>�db]G�Y�Q[�`5hm�eS�h]~�����mRB[Sg��i#�!Ѹ���(X������iD���G��%ʻQ0���:ü�o�'��`���Z���q(�5cH������۵L������e$��Z�k�z(ZE�)� ���L�R�}�q��|�ɺ���4+���F|Yn�PC;��E��X�O_m�i>ù�T��|䧦�ء���.��x�-�n��(�7x�Q�%����*�Q�1�y��x`��}NѾ�A�@�b��E�0{��c�:a�5��љKr�"��q�@�x揬W%@a;Y&{�?�i����-QTWfߟ������I l4�c'i�j��Q���w�������u�溏�����5�*0Jx������$Ke��R�'�Ƥkx�NҚyқ�,�ڈ\�G�F0h_,�������/�P�d�#10j�a1��Mk�3��nZφע����ǰ]�/��5Ch�q����k��va+����k�`;$�.�-���f����9i��R��^������P_�w�V`?v��E9�X�SL���c�fX��
;b���G�r���SG�h�����H�@�Ousަ����pK���#���c��5$i��["����?�g�'l��I�he%���#WH����Ʋ!T�~s��a���pʎp��X(��^h �&��j^��Nj,�#Tc�<כk%�<��>�2����7s1V��@?F��X��T�zaT��h�8nΪl��T�K�!X$�PcȆ��83��ʾ_�j�@�;��(��l*�4���k���2Oi, �E8<T��2Q襘<B�(kj������vg��z���a����1нV��$���( sOH�����]��W!V���������U�(ִ���KK�ҋ�p�cH�V�Fi��z$b:R�b����㓖p���k��U�e�������y<�LtR)(�"�dW�|d��z�A�#݇4<��:�t4{)�nR<�*����#�n1�:ܘ/�iYBl�<�b9%0�aY �/�,��hi��7:�?�y,[Tk3P�DzKsO&ϵXڪ�9�;�.k�P�>�G�T�3+�2�A�^��!��	Y�`3�%Wj9t��|m��u�����S���pC�cqJ��a�R�4��_�x�E��,��Κ��to�����/2�o��jBB���-��
���gI˳����?�����5�]�K��Q����)\�zo,����sذ�����;+��$�r��P�m)�� �lz#��4u\�^t��F
_��F�%OYOJ�H��:F�\I�
H~��:��(�?����4��+�@�j����Z�X�g �ӌ_5^xt�Pno�_�+�`#�4˖�<���8g�����%{N�B�