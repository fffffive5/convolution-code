��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L�� �ٵ�˔�Ω�4�ܛ���7��Ͼ=_m��/ ��������c��i�Ԃ q��0,ry,��`��t�m�Ũ	Fը�uV^�Ծ"���z4�L&�S�
�����c�0�κ�����a9��F��pt[����Q��II@���4�c���a�yS���Ug'����A�U[?a��[�)]�����6���r�i��x��p���P�;��1��$9�*Eռ��g��G���ouq	$=��x6��u��a�R~��g��iT��s��(L4���.�3Q^��=�wD+[�_ٍ%����l	q��W�(�c89�E���
z��*w�$D][�;9��A>�z��9P���T�%_�gq�l�%}uaB;r�Ѭ[v
�{�z6���ƙ��q{Ip���(kJ���v8��4�r��g�"����2+^ݎY#�;�C��+'�l~1�V0i�kuv�䡂!S=z$�p�o��$F��lV>=�t�L��'|a�O���������h�:4��9�1��v4��g�+��֨'�ML��v��D������g���\�H���r�hj�~}Vߋ|J��6ifc�|V��ݔ'K(D�}u�?��'D6�f�Rw�4˸��d9���q�ڢ��/�"�lD���5b5t7�5p���c��#�goH��z´C�t�r";1)�������W�Er<E'��;�-�$y2kK� �h��ݙ�|�鳇��3el�D��S{y�BVY�H��)!<AВ��F����2�|-\ĉ��
S�+��)-���U�5�E`��s��K�X���#*R��t��h��z��VD��{�r
Ⱥoȫ�M)�s}/o��I�k2�R��cx�+0��9�T���Wz���3�@k��������p*�Tt�E�����î[K��!��Ɏ��H��<2�݆d�L��T�U��Px\���)��B���s���a�ō�*P��#'���q�^�F��%*F�m;����Y򈞧E�"|���	��^N�#EQo�o�~t+���R�ƙ�Zo�<�⠃>�|/�֋� �:4P��977,4D樗G���K�w�;�~w���Mni��Ē��q�\�����,�(�5*7&�����{�d��343j��Ӡ�m;⻈��C���X�
6��1����XXK�?#	�c�!_A5�����7�.(�.���PZX�C����#\��_1�?jJh���>Z�<��4���^#tQ�ʓ�<�}���W�5`}�DB�=��\`�@1�(s�A�C�,@*|B��>$wu$�_�f����#9���>�ܚOVFE1)g�-"N�Я�5��6�)��7���:���%��-��G�ry5D��c���ĶI�q��J� ���e���Y��6xsw kX�����L�=BIv�(�͹��K,�Vw��Qh�:[%�*=�ή��#�E��5���c�Ћڀ�Ui�sn6�E2I�z����D:��0�1�p�֣��|O�di�
5z��A.�2D~�1�c��d?����R7̫}�?̠���w
�v�D��Gp�4I�3���3�RoƖڬ!������e_����۴b?cn\� ��Һ7�[	s�;;���itV:4U
͖�x<>p�����C\���it[�"����]���"�Ȯsօ��3T<�.}6�7����B�eo�g�����P.�`몳�[֝ZV9� �[0�Z~ K;�q�l$�s���9166�5����Bo��b���j=��������;g㱀Cv�~��YV��,�u9�_��f^>�QHr�b�X����EuǢ&ٱ�<v�����d���^G6�ʲĘ$�gN=²jE�yЁ��ӑg���2���b�a�iw�|��	�I��T�����-�]v���-��Ztͧ��Y�ܙ,��q�����z�f{��8ˡ��rSd��}��'݁�1��L�h�D�gj��8���C����B����L"��5ɬ�fkvqK$1RV!$5���M�~��c h���g��o+W���p�1��-�ØMTE�V�܄���R\�`���r>��/㤃$DD�ѬI�p��p��3f�k�
���w_��J
H����k��JBet*�%L}�"��B{� y�;��>�7���Q�����oZ�Qބ�D�NY���]�ُ �!�0L��P���*I�gL۪����]�gL"�"��-�Q�-�v��X{is��o�r�}&qGp�t#]K�)�����S }���d��M��+S�a�f�l��KW�yM��Btj{ O�d�&���yвK��(}���&�%E���%>U�S�˽dѬ1ي�6.�����Yro�n����P;��E�"6�{�.7���g^sjF�n�)jF
�����1�*�>�� �,��SNǾ�4�(G��s��#�US�C�]ۿ�k�Y�����e��~LZ�&^��k��E`^^^A��JY.�)��۱�(T6�I��#kgj\�l����1$@F�������aN�K��-��������:\�>��]t�=cZ5�F% ���g�|B�Q��*�8���26�s�ڭٺ�!]���kd|�,��z�Aj�C�_{�Af�T�:ZB�7���,�dI����B�XSe6LJ��%��� r,��x/�z �zY(�㢯6�׻ ��JwS�������B��g�(�f^a�W�"0�X{����)X�?3ȼ��4
���k����T�`����g��ˎ�L��c5�cy��� �IV	�qAN`s(5�u�n%�PSa[�##��QeH-x JrL
��^�	�G�9
o
�L�n%~
״�p��N,-m����0$��!,��'�@�+�1�G�^�� �6�d������&?�v;� 81�-<���*_#ρ�{��h:�����[�YqG��o �j�b4F�Bc�!w�A'u��.�۱�	_�-A�����	9��}���J����@F�t��<���=��:2M6]C�����qN��D�c}~�f%�7S�VN�a�]�
����cw�9�G�=^�ACa"�g����a�З&�u��fp�i�gs�:N�&�\ח]U*�uک�~h�4�}�E6p6G��S�K�~HZ��i���y���Ye�R�S�
�u��ů�&����TY��!���h�J�ݫ%<�u	����#��h$m�����G�(�Y�+�ㆻ+ߑ)��M�W@���d���pG�� �E�3��9�_ɲ����$t�#��?m[����h#�,y��+Uij�Ol�3�)(
@�E	�i�V�(��U"������0���Ta�@
p����G���$"պ���Q��#8�G�U���Wŧ5������d�\�[%g��ӓ�%�J}]8Pz똊-T�2a)��>I3J�A;�:\p2��QИ�a|�r��$ubأ�#4/#���ۚ�!�g�%�K�[���wE�R�3=�4��N�>�ҵQ�q:U����#������>�%|���}��
B�u��Lm��=����$1�b���s��w�p7t�v�G���1�
ܰǼ;��ɟ;�һ�b��~}�7D2�� ��� ��c�C{��R�/e�[�]�af���=#�?+3��@R��3��y��6 ��kzQ�iyR�������[���a91:˭< �2.?�5�[�4l�lY��W�0	Y�nz�צȥm�x���Pg��z��?��:J��O�����N�o#tRhJ�:��Q�D�T�+�i.��D!Rܧp�|^�����!�}�ii��DK����J�ô������
f��(3�2�'�C��|�[w�k����Sy�?�ݣ/wO�ؔB�0X;�~�CD�c��Nx;U�^-�~����f�m�M9h�@����e�Z)��E����H( t��6�܋����Ï�c}h����\m������^�P&�C�TUy�%� Qq���U� 6�����һ��,��DmX_I �V�0� �� i�C|����ߧ�hvY���Y�q#�Q�?-b6P�le}���ܭ��W)��>���^E5{��$��g�|gj�P���aCl�2?a��%�]S�h� ����9*/-�ٲ��F"���������5oWll��+�9s��ޚv$R��߃�*@m+c8Z��	>�Pc�L����I�m�d��s�9�T�)ڰF��P3r����k��Q=d���1Q�).�el������\箾�Ԃ��+/�j���|8�j)4�X�� �Ʊ��vx�s���Fu�Z��%�#���F�ǌ��h��K�B}�:�%#mA�s�}�%�m>B�_/�$NZs�Q����'�AA���!�������^L>7>�GPNEhkZ���<�\蟎[�޿e ��zi�	���ׯ!���ݛ�k�R���W#�K4��t�e��=D��nd��-Cp��d��PAC��`Ua�K�&H�م��f�&��J>M�GUD�qy�BXB�i��]�q0:�����Z9/�/����6<<��;�]�Ȩ塋���S�Γ�s޿  �h ^�w4��"�����v>nċ�VD�#s�˓+�������\ך��o�J��b��Qz6���	����A,ӄKȝLD�z��@�27�3=UFk��7Y�]{�D	l�m�S�#���� �[�;K	G�n��nNg�zz����9`6�V^w(Ή�}�ؚM��a��n������$�`pQ-�Õ�3��/k�id��&��o"������Y�<m^u٢B�q�H��J����pWT`���[�f��@㝛�@�����;,A�ʟE�Do�!f���G�T��T9���Z�/�z��2?g���f�J'�7AЉ�PV,)���	���䤆�Ԉ\Q
���W&�x�+3�W �����y8z_�������� �|�K%�s���JymZ??����� o���G�w��V^V4|w��"�t��\�ֵH�Ս5��Z�ܑ�k�z�"0��y#W����W썎��;CF�{κH�#�4�����x�(ukx"^~KV?�r�^��#VXֵz2L�dARI Cv=�k`o��Z�cX��r��@�'}-�j	�OD'J��G\P|i^}�+�[0��(�x���V�M@�L��N�T&�3���AÕ�-�b� =�gl;�${��+�~L��Sß�Y��N�����Ӽ����i��g�e�N�)���MV>X�)`����pəj%d`y����q��DCߊ���e
[ռ�V��w��y��1���e��;A���Ģ��e�i�Wbg���wNp)�y���Oz�?9�iڅ�׃����l�3��/���P^�C�e*X ����r�?�cנ ԁ�5Oz�L�X�q��c�mȾ�!ij��Y!�x���޻�t2#e�ϨM ��I�`�G�h�,�}��h|p�l���>�(VY34���Vb��޺(�x��� �3l���X�"�-d����6����O?_�s%�&��'�:�:X%%�vm���7x����h��9��`W�b�B�[��IoM�K] �k�#��>W����KM��E��Η�t�F��o�6��
�K�O2��*�z�a�?�l�$ڈ��W����Hd��VN�u�Y�J7���Ƶ?�O�1�Ӥ�2�>�
�W� ��|�ct��1�ݯ�\ho��:I,2�l\� �䲓������}�7�t��&�s��S��>0*������pي`wD^�R�9xL��t��2�������=粒��n@|�-�<���	`�^�|p�%�~9u$#����J�-��M5������n��5y�x�3�vh����w�AA����pP!V1�*�\󺈔�S5y��Km��顷�%�N���~!D	�ծC{�pIu^� L��������.	���8D����r�®]8g��LƢY�TK�� ���c���-aҪ���Ξ�:��������ƺ�;��E<��ծH�u|J#A*R��f�A�����h��7��{&�^ꈵ�Ӟ7��*�z0nP�l�њ��It���E���0�;�e��b��>�)�z x7d�G����lxwQ\pST`��bK+Q�qA(�y ��P?�-�Ў�'MO�L�m�ϒ��c�ui���Bf-��r�E*Бᕪ��FbQ �:�DƟ,u��X��Z�_���p�?o�3�CX9���T�����Cȩ.�G2�7)O���+ݖ"\'�R���3U�w�����,�������v|��(2ݥ�zZ�� ����l
�6��@�0�)����z7c��J��L�hH�%���gj-ҍ�0B��s��2뭇�}�oaT6�;8H�CÕ�M�M�U�NbB��u �p=��b�X�e���!�������&lf��ٿGĊ�a�4��)��X���s8^��U��%$����XX�GBf��K�g	�G��D��z��0��	��H$:#�?�E�ܚ$H��r�mQ��V�<8�H=H��S�������ѢvojД=������Әʣ�Q�Kk�/n�b/ ^~_��9�r`TƩn�
�@-��-wC[(�!��C���<N���૙g�آ�sM-���;PȽ*f;�ш=��R"� 0[�8�x�}u?t>�I��q,��aR��:�����9J�)��fe $���߿a��K��Ae�5�B���2�:�|qT��Z�	�`V�F���kj��+����2��-�.sx:^#]Ѱ҅<(#*��IЏ��Hnj	�"]��.�{��U7S�͞��=�}�uG�Mx�"�n��j������������Jm.�＊�$�u��4F�06���d)o���[߻��PǮDa�/���zP9�=����$ً �����iy:�63$�UJk��22F��P4U�&Ł͓_k����F�vz��r>P�ŬEv	��G��JW�o��G�D���_>	m
q�:�**�R�Ҡ_�ʃ攚�d�M&���VB��>�^3�<�$6gU�+�c��?�bU��q����������'w�j�E�
�D�z�Z��(d*�<��>��[��T�"b��7��j��3<\��"R��i.Uw��0hG��̐Z+j��?�G��/�Pc�=�)O��Y�숟- 5�N�"���h�۽�V
�+j�U�ȿ����1���$�K�H[AZR��guzi�>__�-,e�|<��.�EV�J���;�I��F��c���7KT��������azr�*����!O��DK���Y
v-���k �������H}�v����4�h��W����~���}n���*���ژV#���S�ߍrB��T6�J��P����ɴ���{Р�Md��rj�վ1�a�SM4cz��Z��Ur �3�P�����8�bl^H#j��-!��M#��M�x6�Uz\B
J��Ҥ\�Q��&�,+��&�Ҥ,�'��������cֹx�m��=�b�dː�(���Xu��c�/s0}�z�~_�a].l��lӜ@Ɔ����N��iK��j�|,��@�y�<�}�(�'k�H��� }wcU�[�l���S�L�ce7Ŵ�-��n��m�v�!ݮWs��p�њ���TK�c{���J�^8�C8˶[}��b��\�F���-��e�z�:�͏*���u�3g9�:�!��ҋA��*�y�+�i� C'G�@ቕ�e�ԷFV�{ɉ媗�<os*I+��75L]�f��}`�gb�V�O��dǡ�	)LIj�I�L��F�48?:A5v�=MA��[Ih���C�,!�2+�ڷ�Y�@�$Ҝ�k?U9���M�8�y�7�K�)hl�D�) 4��[��/��ĉo��T�]����s��m]��g���(�I��-���睸��|9�In���(���H����u@�iN ��Ҿn�L��R5�8�o��vd �6I�aV�"��ݬ��Fft]cfL��%)P�ԁ�l9��#�����vp/��"�Kj6�R���e�,��P�6fX���eK��ݺ���F�r��a�e���X���� k���q
����8/ WJY.d !e�+3��x�i�m!Hâ�G	>�ʻ�@蕏c9�λ����Ě߯�7��� ���ևb�΄��v���9�-��1%���ptvΟ��������#�I8ޭ�"�G���
;N�q�Gݞ�����2��zv.t��E�J�3�3�R0�q̊!����ʄF����z�(lI���י��f�BU�#Ȁ����ߝm�o����H��,����Ej�p���Z"��؅A/�C�z�J�s�_cl�������-���4��|�9�bv��}I��B�)ݓ����R����7�4�A�笉 ��ۈ�-3�%��I�mE�96�[�Rջ���ٸ�͂69-RC���{a��}��+l�2�S�H:*n�
�����b�7��$g^v4I�#TԳU���íz����� �M��,�zm1�S����"�ݿ�e��*���o��ެ^p�<�S�OÌ�e#�Q��{�K�F�?qLk;��SV���*'*��n ${o�*�ژ� �|�c�1����w����-���{��GXAR��/)�������	�v�N��?Ue0��pFB��I��n�E�pǟ���
���̈ H�@]�h�י��8<F�[������"˲$�Kn����EV��ͥ�}�9[�~{��*D`o�}�[��|Å6pͲ��R����5�*�*��n#:����W
ǹn-�fZ?��z�./�i��q@c��	S�"V�#�\Ij�w��@:��ee)cꡲT�(V<�QEE���&ϣ5R�x��`�d�f�V��X�v�_���6n4�����r�=PnO?�VS�C�?�r�q��	��"4����!sq��\}B����Oz~M��s���v ����;ֹwg�dv&��Ş�\�:}��K��q>f����"��b@d�4�+{}2��E{?0n���`l=�η:�Z�-��
9�B���s3����^tx�h���:*���5�UC�������`�Ze�:��:>� }�<L<է������|2�Ө���m�o�O�w��	�Y�0�Z���x)���
��Cs���tTr�krie����sQo�/G7��L�Ɇ�tr$9�ן�Q[ʍi� �#r���ۖdh�4K�`�߅����Q�䴄w�yy��W��Cg�>����GK @T{ێC1��NFd�0�h��w�X��`�x���.���Ǔ�oh��a���&t�?־HX�z.�R�
���D��5ҷ;IJX�K.D;m*	���o	ꖢ�Ţ�C��H�Ȕi,���H+�0ˊ+ށ�y�\n�j���*���$��}{s��O.�bqN[�>s8�p��8�?����W�MJk(�2i!O"�Z��&V��1|#��8FNv;����m�\ئ��[Q���4N�Sz�����g��c��^p����9\�u�z�Pq$L���[e[E�tʿ������͙b��[j�:�0X�=ƞ�bG-�S�gm�H�@���t��q�4ʜ�z�S��.7G�K�P"A�S�0�i��i̚�ɸ6"���*{c߶8`��Yb�e�ʍ=f�k�xn�m�_;��b;�������ᥑP��c��@Z.<�q���3��4�Hh1�7Z5�t�X1��'V�Q
DQl�V�9��akC���-j3XIgec�WG�T�Ozq�y��D7�zW/D\���峮E�yi�=�����b?�J�&OB՟<=ꗩ6�X����O�Dŏ�!N�0F6����"F8�K ��Gɇ!Pm��л�E����r���w��0��16��G#}l�����0�}�w�4�����t�1�,�nC�˻p��p�����#��+���$I,{ES�b����/�C�!�$,K�f��Dn�u�Mث�@��5���H�(�Vg��e��J��_�**o�Pj-ny\�]9���FГ��
��^�c��l3�\�����������U��ƠV{Aܝr��h���V�(U�Gc��Ǥup�SW枉����\ �j9&#R� L�I�C-"�.'Bk�@Wl@�TY<��~�6�20�RI�6�����x��<�uD���F�8��0SJ�� ��v� v���(Eg���2��pe��\<�ӧ� 	�S��퇗�k���G�:��F�D��f�w~�ꪲZL5H��iz�Nr�|s8���(~�	k\I�s���`�3�3qjm�4o|�W"�rE ��׎6��}t'9)~��6v�	�tܦOx	�g���U��ج�ҳ����S�9���A��4�%��A�qa�3QY��0��1�{~A�j'T�0݋�;I+�i��oks��M�� �e�[0?>|~CHv���%��Y�`�M{Qo�*"]��pp@E����RGȴN��%�h/[��~��宀��_C�.��@��f�|�)�wk�������A��e�#�-�}����<c�Mi �Ƈ)�%��J_|��0��=�\u-=��%s�u<�jA>��$�C���Z�t�,��Bc�{ic��rg�;�@]DY$��-C�����EDdH�[����H"�iz�n'�);�=�u#�s�d��i FxK���a�%W<{Ǡ�/=ɍkE��lh�~E�	�?�xU����g��
��Z�-��"��T�����˯A����ƀ��]��ٗδ	~��
�c{:F����Y�,_U�,��M?^<�h�?��v'	Ք2A���Z
�rg�
�jd�g����o�%q��in��iU�����Cֹ�r�c���Dy��z��#2<2�l67�x�E��`;;�8�x�T�S!�:)�N���鷓���;).����:�����z2jk�qK��8�l�L�+��,�P�h���9�m��)�i��S�)ƕ�A�g��3��e����T����X����'|�꜈NS�����ٓ�i)�Ge9�t� P�4h�9AxG Z��Za?6W]ePOV)@V�'�߮r�Ja�y�0�TKHΌJHLsA��2!'��R�<|�H� H��#Mt��� �(�W!�w2xaD?M��%	R}k]>�]|%N?y��Tw��-���h�,v�#Nf��Ai�y�"��������ȥ�YS>oj��T�Z��R>��^A�zp�����Ӆ��S��o���BC���}�Ę6N�Iʜ��1T�&�0S1b��̑`�ZҀ5�C������L�A��);Ν�V�� `����$t�Rm�~��[p���"���^F�FE��
�bsV_���E�ޖ���Kg�t��W�-�E�(�����v�C>"4�"�ʫ��Y��y�i(��ѳ��t�5��Ċ;f�mA�X�H�δb@F���Z�~���0�iy�ɇfs 1���|CP�����O��y���6�z1���L)]i$F���$�2��Pc��OK4��/��(���V���<��9*&���,�g7o4�z��?�@�Wޜ1�� ���r��vB��';�t�#��<_�R�.{�,��+?���gbL��`N��35&�ⵍ�¨�H߭�F�|����L����e,�:�Y�G�"v��$��$ӿ����u�x��ՈN��C��he�ȼ��B����?ce^�$I���Z��FJ�i��/��+���o�+�w�M�IQ)�! Qg*��T@n����
X�2�ܰU�&T���BL�}Q�aBPk*%T���@>���H/˅㔥�����%�v��������#��|'��ޛC+��(�R���xDC�����2��Q�&k�E���N��7©q 3qweӃ�ޗ�ҿQN�4�5bh��C_4���'��"�Q`�*�`Q�D���|p�����[�g�� ���������o��hU�'0� �V����K��$j(=r���?�/�F����EQVI�>���p\�H�O���8���d)�B1G\uQ�v��]ra#z.�\��j��c���>l ��n�`����)-$���r�!��s�ɍqЇE�nH���U�w��$�lu>Ԍ�˻��i$�<ڧ��u<�q"��v-5�*B x�������q��D���/���\�>Yyb[���FK�V���북&ׄ�B&@����LYt�������
-�;�6�j8/S�Ԉ2p,O��C�tWm�Ջ��Ղ���$pf���l���������]��Q�5���/]�AQ���#���R�*<nm�u/���/�c�rPw��|e�Q���O�ɂ����y�3����V�:��f��Rƿ*]�/�a=��c
r�8��������\����k��<^��~�qlU1�]9�QI�����Ԩ{+M[�z,�k�Pַ�>|V���\M�ā��7��P=���3���V"�7)0�L�IE�9�6�P<��K��|)O��l91�|��N:n�sW��,�D����|���}�[�K�8�Fɇ��r~�ڸ��=1�`m�����N�J�潈U�%؉y���U���o��KϷJI�2��WeB�@;�D�7����s�������o�Մ��y�=a�����Ҏ8��i4p�:G���9T/?\Y�^^���!�uhz����B��Y��L)��Q68-�ďR]��l)�]f?y�b�2�'�ݚ����}얫��2�R"gw�2H�wv����1�,U�;&�A���ѨnprN�m�%���uƓ*��P�YEq�Õe�US�� ���c�ȼ1Y��LC�r�Om��A ;	r����l��+�g��������ΐ�l��æz?8��Ooe�j�*��8��0SA�柍��]����S�)��϶��N
��wgN�WH|��%�?I��JU�^.ģ��I�2��I�/i�[�1�-�F�wH�k����6���Fp�)�v����k젠3���	W�����C|���Y�X\�d4:�q�˰�O��V��'�p���Bf�`���1������ȧ	�����4}�MJ�5�r��S1�קg%�>�9?fc`��e�w�~e��t���C��'�=�Y�����l$eE��[H�+�4\4�U�X?�4�\�D�@
�9� �L7�v0�%) �
�ۛG�"C��IP��ʤߠ����������*����a�ݸ�\��;ֈ*������ܙ���jv��V��/8��+Z��\�4�jP�o9�� -�Y��V>vU��`�0a$���(�v#�aY��}#(�2J�on����#�/1j�����U�r�y�s\O 	�����^jE�U���e]3�T� �������6_r�ız[����F�جUo_�&D{��Y����	��	/��\�j˕;`DY*�){LGh���35��ki 7G������5y����?8�G���"U+5E��_)=X��#�=�_�߁'󹏾M�f�6��,ɝ�����Ш{=�Ŏ�{$���@Z�x���c��h�ޗS����k(���ŝ

8��@$oǡ��r6�E���.~�Y��� ��Z��Aƭ♵f-?鴳c*��@i+���!��ʆ�������Hɦ��ǁU�}#�'�svҵ�p���'�Ž��v��s(�g�T������o���ҰYX Oن�L�!β��83m⼐��X}Ҋ��#�GYm�97�=Fiks=nNܟ.qJNfms��4*^pĶg{7@�W��.���k���bcյ��i�=�\�}�����&�E0�%f{f�[�N"a������
:�j���
�Mj+c8���J� �%�p�@��;��;�����>� ��ϊO���E��&��U��F_�:��eyUH�3C}^��.О�*	�gM��F����-���?����Ph�J��RZ�H�Y��.����O=�����,�����gUHZ�^?��i�'p\�/t�`�*��i�d�y�'�ޔ�����ړ�)��Z�^�=dp���9m��0F�ۿ��0�n���:������=�l�EZy���sd{����7��Ub�Ə��𵋘��j�e��,�^䛎zbf��|�Rt�a>���i�À=�J�Pr�I�P��Z��!�P�����A�7��?T9/k�d+��Ay*�ث]�À3�=�0,�Z-��Z���P	�s��+��$�%,ξJ<� :�~klp|�~����3p�Vj��������V�/&V�{�(9�amm��/ĝ��C|�*�s^�� h��M�4� ��	%eQ�z�j��V)ż�PO�����5<�t��,��'6��Ǜ:K��	���@O9W�����{!�ʝ͵zH�\�ӷ�Vⵈz��	��&	�g��ǰE���v��V�ت�"A]���jPP`c�����D0�
�8'O��>�ۃ�kתm��{0J��E���j]5�3ղ���Y�BƘ@�0�swf7'�D��41�Y��ڹ(٘�'k�.:���F\�&����D�qFV�2�U���(k���=��eL~����0&��C�M�kH�� XKͨ�)-cB��e�Lz�y&j�� �����̕����٭ke�3�}~�S/� ��!��U�;s+rN�.6x�X��Ey�F��Æ�#^��YV�>n���2]��G�u�ѯAsd���^#�4���l[��A1q�$�W�
s��	ϰ������o>SͰ��E~���ڥ���ͥ/ϞD{:����������/�~h����=��Z�K?����On$��{���V��g��QgS���&F�nd�)�ھ�	Į\1P~�g�&�X�nm����;�2F	�c��0i�1��i�Yߛb	��a��HX)��N��͗���/8NZܿZ8]�SE �KWi�e�O�Rh�nN9��㫰=.o i�y�H�Yx[q���_j�N<5�C��RR����eο`Q�R�T������:��jIĔ6�ts�5�xh3YZ��6�s�W����N6��W���� ��;`wa�zT�Ќ��1���JW�c�ȿ�ez�� ��ó�po͢r6��XB���&�k=�h�X�1�"v���T�����|�pUhbq�.Ybń�W��y8�Z��*�jD��Z�Y��z����g�lt9\"M���.y��D_,7�ܶ�S;A(!Jy,.h,���E�1κ����\��BS�S�~��n���2�J���'C��)�i#<i �N"u�̺̜Tp�ےm�a �AJ��'�H
J�D>:��#�P��ؑ?n-�"�n�5�@'X�G�S|�A��	�kHO\��յ�� b����{a�oJ��?��ڠ�	\�;VD�A%j���@δ+~=,:��A��Wz�$���zo���׌�w����F���!�[����o��	,: ��I�����oPMX�K� f�a���c(:)�~��M���>����c6!�W�7�/�Y,.Ǫ���8IiLP&���7��
\���\���\6�h��nǏ雮��u�1P+J�T�L�LVn��	˻LB���^���35�z+��礈v���(�(�3���aʑ�3�$��h���ksq��_e��_�c�	�W%����g�T�{�R�W�>*-����!���O"���Ρ��ո�|��a�yű)���mQ�Iu\�ѝ��������iל(��[�����������UW�N7M.�L�u�]#m.��Dތ�6�tX08��E�`|-��@iW�f��A��@%��is'�:丂������;6<�l5����K�F����]�!<�O�$дh[>�Bߠ8�D��ķ�<�U��&����5�,{G���0482ʕ<��������M�;��T�=������x1�Wn�W3$ϥl8C�wtɻ��L��L2��D��`� qN�zNˢ�/��"��̏��~�lp��ܑ�52��v<�b�⃖1E��zcB����α��6��k����J����g"���a�$�0y�N"18Z[�%�嶘�(%��Oy��{Ão 98�iT8�3Kܰ1^�~|@/���C��`+��=š��	��&�WP=]+����'p�L��Vj"��a�3�py�0h�n�#&e�`�6c��0bvM��+$ڨ�Yw
����+�C)T�p�T����g�ޫ�F� �5�H��g<5��^�& ���0��K�:��\66�JeC]o� �"="���c�"U�ҦF8h���\�V�.�+��ʗ7f��f�W��ڃ�2�B��@�ERD�P�|}tSP��UDv|;�Q�ݮ��h��)����4�N/t3�e�/xu��<��ySp�ڕ �f�&>?M3����Ca8�tz<�b�1rmú$i�] 0>Z�-��L��8��~N�o��CP$�
�<0a!�r����[�?-t���;�{@-�h����D����i$I6����ϼ�|u�A����8�w�8��ה��q�*W�B��� �ZQ�cb�$�Fc����<kq��Q�����a�pLEX
�h���yd� 7����=��}���\�f(m� ~#��g�4P��!�k/+R�Yl��Ն�:ȭ�3G��
e��W(W%���2��1�Pڰ�AV��p)wdkО#�7��V�YT�����h�hW�Rܨ���J�_�q��/�ש&��v�́{�����.��1�K��D����k�i/e�d�����E8F�)�qH����ފ��a�����m3b��g��ڶ8���G��U��^4P�t��5N����]��Őw��$�����Ȧ��M�{�
kLV'm,2y �� ��n�;�.a��Y��`20Ί��thnC�!�q�k�x ��Q�c�}91ld�´�vɏq�Nh��N!�-��&=al˝k(����S�T��_,��*v��"�P��C�����~i<�A�WY�u{��hڄ�N<`�͋J�v��GiDߧ
7hw��Y��7�(�����1���0i�aOy�} t ��cAN���S���f?B��@e����S9�~�����C�d?jCz�(��ou1e�hv��~_'��e{aKD8�~r�/���z�Aʵ����'b,��0$}�[�e�Ka�9^HՈl��e@��"7��y�8e>�Q��qn�G�tƸ��� _%�t��RM��N{]��P�! �= 7��'o�=�Qi�N�S.�z�kc�
@��ӭY]��M�[�
N��'���"�ͅn>�v��d7�7@���Y� u����,{��*���	�}1�]k�9M5@���=[�n߉CR�+<�c�Ԧ�OW���,��tNNO39�gs��Z���Ml&�ᐲ��؉׋ 3#Wa�t=,��>���:O�f��|��i9}Jzq��M���w����S
.2�J���q�m�OֈO�Z�z��i��N_�eD�].t�0O��۬�$9uJ[Ƨ�)1oql�^W�^(˞*�- �a�?*�r!��@�&݂Ǆ��»���CHU�a����<�eT���.Tؠw�oף��M��{��0���"�����-�j^2�˽*/�yy3��&QNQJ�:�=��a+���i�Bֺ���8��(�Vd.�"O��]h�8��0Y+��h�f�
�~�`e��Ms��y�x����A�7�������[WQ�7xH�ی8���7��B�/'�Ѧ�6,i��S�������p�ޗ_���kq��y
i�����R�(�؉.�Q��#=�KȢ���[n���t{~���E6�3�s\)Zg��G,!@�T�3���W��\>k^�_"���6�>�D��$�$6~ɫ3��/���o�������.Q��#�p���恞���"����W�����I��<�����3k8��rkr;-�ΜR=�&���on�7��wǀ�sb��붘�A<����:�߳���P�3�y�9T��;�T�!bs��k�h�����)�7|��rSu'n��J
T���s�M4`5}"�����#d�/x�N;�!�1������P�L+�Sπ(�	���t�MU���n��|�4P6�V�O�*�"�3%�%k����z<�+Gq���X9���k	L�����
m�c(q0RNUNw���g�.�P<��þ����"�L)���ƥw���݅�2y=v�1B�ցߕ�U�y�\���3�Eqh�����:G˜]�A`ln���k��̠80�!P��ۓ������&�{��5��.�tM��6x%��z�k"�5�@o7`��zFح$b�CD��>"O<�`������B�J�l`O%����Ӓ��7փH<�U2������	~3��}9P����{=r�v�[���6�NmBg�.���jI���p����Hl^�ӛ|�m��=ð����wik�,9�jF~ڧ��S*���8Q�rE��t�*%���qi�oM�V������w� X�SV�z�g�d�+��W���U_����[�@�(��/\��YX��.�?�混�q�/��Sg��x?6���!k���I��uqoBLz�>����^�s�#b�ƚx�mڝ�Ԙ6���xk��sM�X�����Y�����հe=��KY�Kq퍸�"�Q��A��b"5
��,�ֽ1Ň���ыH�2���\[��^��:�Q��㮫��o(�n� �xd\}�,��f��3�r��3��M��*�7J���wP�J���X����.�'��8ggu��K��]�p���_aX~��;�gNJQ�6�G�<�(ҿ�8���v�򴢋�X<0�GIى���U���2�lv� �O�g|�"_�^^y��i�|S_+C���a�q\b��}d�(	P����3�aMa������R������V����p]pR�ņ
 b
z��
^���5��P2�+%��1��YN�1.1Y�l���W��:c������w��EO�j*���ԮE�~��ʱ]���N(��l����������"��MO��O��pO��ACB�1�u�g������/�z����?�Bw����I�mS��M�ϛ6�:��t{ijw�f`l�62W&��7<������%�l��.e��/�I�_��q0��6��	tf���m>�,��Q��-av/�z�M���7v�����C�r�=�������jRzl�ee�����01>�¬'�X�g��OE������J�1�,_BPݫ���)��b�S��[��ٛ��d=h����\@�r��(��{�x�xE��	��2J�E�Y#F
�^�#��Z�pm~7ٕȦ<KO�r�И|b�Q���P6g	�	�]��d��9L��{t�ဆ��lǵ�����]�(��E������l��Fq�9����U�-�U����>��$E��>;�3�X<�'�+�>�R�#]x��/��*��[�X��$w���4��!ދK�� �uH$�d[6s�����s-��<m`��Wf����z�BOx�A���j��ԗ[�&E���}�oV�<�هKD@v?Q�km�0V��ǀ���Z>������������ט��O(q���Ձ�����T����&8�X�~�r��.�Qd�ʶ��&�w��z�p�v��^Aб��`���l8�^c�T�!m��z$�"�'��� Wx���3������$������w�C	sT�x���8��B�Tӵ���j���z�5�b�SV����{ػ��\gm����2��c��B����N��oY��wvG����7c���n���_�S����g���6�'K1F�E�g+�v�.��Vύ��L(�T�"c�qC�M��@��#��MT��܏�����T�/.o�Ŋ�ֱ��� �����8��+��._B6M���.�l�]�cG��B����.��qX�.s�������-E�o���t��5��dm�����K>S^����H�h�U�0�\=~^��ʧ3|7u�c�TQ�x'�(�3*O�Ry9큗¬��8������#�~b�y��Aپ��ń��>��4�H۰��2�����G�0b����1v�N�syv����c/���6�ssq���D� d��jX_B���)u��rFV�L�!g��=`�QdzmTY�DU]�����.�_8�/�̚�_��ٔ �rD�U���ܐɗ��2A�$"��I����i��~ʺ�>�w�L8�L�Qr���\���t�1��sf4��n�q��N��h�����O����Ϻi/�QV��S̱��!�_�pە��.Մ�L���q���q���̗��B�n�9 c�F피oO[^��0���(�$VP2�B��"��Fr�{�[k|hl��n(Y�u�)�E�3�g�U�uQ��D\Ol�^z]7ˎ���F�2�խ�A�h��|
�1&a��=�uٌZ}���:�숪��s�ӎ��6�o*|M,��d^Z��w[�	3�Ac��<҈�����ʻ��M�fT2<S!xⴿ������S�o�U�E��YZc��.-�r�	������F���B����3��W��SAD4����ɨ��@��y�5C��+2}�}�y̹�je�M�)���Fk"��)�4���i��9zu�9�U��>bu�����0��?��n�Q|�NX��hҮ҈��n 猦�1hx#W_O��h`;����kIns�$��K|��� �l"e$H�gh2�����.�C���'62�
�Q��z�I�t�hf���"��\F8��"@���o�Z��֯B�1�zx(��Iy`VK~�ˢ=�O�m)����u�ܷ	��:(|�ѳ+QS��E����j�X���h�ň�?��щ!&����q���ׅ��4��;�kG���A�
��k��#�y��n~�t�����+I���}�o���8ԋ������i�4�����4	��œ9�c��!�Ԕ�Wx���6,:�i���q���J�$�D����,���y� ן�$B�r�oL4�<�h�M�g�K�#x����i4ĴD<