library verilog;
use verilog.vl_types.all;
entity Conv_code_tb is
end Conv_code_tb;
