��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<���t��ejk��v�C</T?}V�E(����L����5!ҝ�wm�!��޳��(]$�l;F�$�тJ��̼�ҫ�j�y�2���r�R���(��Z:φU��q�P�,�)ЄWKh�{�~�[�wv��M��$��*�nq?WHY?���6���@Oۡ���4]ʆ�n��ʗ[S�����JF�e��T���%��� �j~��4�N��(L�Ng�O��#�����#t�1��l�����G��Z=6-�*���j@eʰ"���X��������}-�c��F�L��ob�;wޢ���m���f(�M��MBq���|9{y#�D�[��Ϡ���u���$�0u%�6�-�>B׋W�>���sT8
k
A�:{���t��v�qNV�Q=( "�?U�L#�� aH6�X�[���P�
&G��lA%j�r�w�1u*0���g/���zPÃY��d\��;�mCX3?^��M��=c����kc��az�-�(�jӴ:�TD��P5^�Ɣ����~>�l������[:��v-`���)a�RDJWv`�X��ZA��_t�!y=*�E�%�Ex�+,�&.d�����G��G��̏b���7�3|ׇȮ�!'�)
U���pZ`(�S�Cy%�Z�U"y�&�c;'��y�4�S6+#޺>�{H�*���r�IFaFC�����}@���,���_<�~ #�
L�+��nm#��C����+{֟���K����K�@��9��.$�S]��cMaL�B���c���s��"k��E��'P��ȯ�\e�˾�f޲��V'���W�����g����F[�s���YV|�!��="�0>\Ur;t>��&��ǗgSRZ
���Z�o�RA���K��[��������,�+k%������6z5Դ�ĎИ�R|�x1ZY�Lz")@�}���r�`�����lK�F"�����U(�#�'��R�3�,���WzV?l! ��b\h����-�ċ73IE,�����)�]�W�3w�HOT��WC��r2Xh��y�s�����vc����vңD���������2[�1�A�6"�#��V�;_}a����TG����P�,ɲ�*�n6
f�u��%/n��EK�JB�m^�n���I��9� �Ϳ85���®h��V�����;ČL2<�;�	6�����O���T'�{*�B W�q��"*�o��'j;L>h�ڿ:��\D�΄YZ�E|�ԕ�,t0i��=�T�����U�B� ����hB�,h��٣z���3�9���t,3]���&x��w����;e�5V�t	��/ͤB�������<]b���ő`�4�c���s?��6�����ɞ~�D�*�;�2�ik\��XzY���4m�A�,	%�
����\FM_��*�����
��78�|�<�e�X��m���m�
?�3%R��3Ap�\��ЂV�����fw��L}�����q���+ �t����}��u��骉 D��e4�૝�Tt.ւ:�hI�<9}�?�v�<���e[�R�-z݄N���YG��݂�cf�X��ӆ�H%�}@��].��OqV�_�I����n�����������4�f��W6�A!eE���a#�"�)R���1��	�;� 	��R�:L�����_%C���n���m�%��+o�����$1���aeƞ���=IMƩf���l,;��Ǣ��	�.����[�'�5���@֘$:�c�Ag3�M��`Ĭ��7�������Rm-��x��%���Vi�$ƺ�
~���ni�V��	s�9A&TX�A���aU�/~=Җ�zl��@m�&i���lpe��Q�I����T|�a.�P�#P{r^]P�2���=�7�U,~Ps8bA�Q��2^U֤���]$�l�w������S���M