��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L���VFjU���_+ �:�f���E��$7�'��;P�2K�9 ���s�D{�?1� �7�("+M��U
(���h�gқ\ �cy�aIzD�u��B���9�E�8Bg���/��_�D��3k�d��_��T�)�Xzk�٦
l"��Kq襏d6���r�O��+~�����wB�|��K�D��*r��̬U���c�ӏ�ӥ�yZV��s��V�7��W)cH,?���NJU�_+�����x/����0]d�!�����|�!�V�w��'#��g��J�7�]i���H�G�ڷ1)�2����N몏hG
�@���d�p�Ú1J���A#������_O�I*d�}���M��ʹ[�7]3�?�'r�fſ�$���"ZGkZ�0LG�������e�j��}�As�������4#BI��)�5��uU�/2�� ���>B�p��t|M��!2jH�����iɁ�q�0����h�^��lJv��D<<��ᆕ۳Xb��q��͈4���)���c�o�� m8����ST��jiC-e[3�sW˖�{{<��uS���F���E-��+�1�P������í��h��B��1R���P[~�Tƭ�@@o��D�!����f����Հ4�DV���-��R�O�:Y�F�N�$e=���É���F�"�9ۊ��o�-<@��b(d!rU���R�JF����R(�i�Ifzȴ��w�=�]3|�<�T�NQ{X�6���s�n$h�3��O�C�&�{r�=~�O	\��o3�~� ���%q9� ���bZ��q�$ 5g�O=�N JH[�����*�RKW"J�]�Z�N��w�
�}9���P\�_��[0 �7�n��]vB����3�>�a�h��n�k������J��!z�qS ql����E�8Ԟ�K��B�Ŏ��Y��%��a���&�t��+�B~~D�ie3�t�i�:X/w�c�X��.<-I��vy��g[��F�C�Z����h
y�N�3�ʛ%�KT
���7�<~%:��J�01)/m�6)���Z��K��� �~R��o��H���+�ܓ�6�6ܽw�g^L,�� q�w �&4��ں*NNR���-���U�:�n����Uc�7`%�Xݹ�w�;a���׸�����]Y� ;��VX�-��*PEj�����p��U���Y����ً�����"¿�t�:�h`�@��R5��J�?�&�ee"���Bڝ���ӌ��Ё�f�K���V���B�� ��qt./�0���`�)�v��<�2��E�c�u5m�*�>�AޑH��^3��ᾬ��&��T��\�q�����g:�s�v�&5U\tyi9��.$f����23��V+����]JJ�^7.p+5������@���8�}����oF@� /�q��>�d�≥F���"���9qT�;�L���گXF�J�:ؚ��(��(��1JO�"Q zǰ^�a3O#�!���A@�+�V\[�/����1���)��^�iYq=H|�20n^w�Ch�_���,��;�c�=��|�'1PeGfX#x�u�6���F��ЭC�g�����-�@�62��0cL��p%��]��(����2j�8�H�9����OK��f�����ܮ�����~H�mcհ����E�\�����My�:��F�B�ԅZe֣S�c_��f��4��GnH]B�^9��B�(
�o�8�>�Ha�R���LЈ�u\Z�����8֨����`	ͥTΞ�Z�:Fӭ�o}�Ar����3�Ӂ~9!^y�b��Tv�	�T*���˾��D�tJ� S/�Pg�H,��n'_q�n�>����=H��\� p �o(8����+\SU$�̳r�e�C�|�Ƒ���CK��en:�-�YTe�T?M�~w�rR�rv���1��~a$��kS�
$ػ�c�N*+gh9m%8���EUu޸��ˊx�$u.8�d��aW�v�UH�됸1B����|
�WR���H]A����Ѣs�tH�?)��V��G��H�V)cĸ����=(ϋ/�������a������9�W���SF�ӿLl�=]�,jh�ʶ���^p(`Im�X"J̌Q�r� ��i�=19mr;F�3!SRX����]��8j-�a2�^�
&z�>��<��|����!ȑ�_�v��͒�?�jQ��4�fA�v�� ���Q�b��j��S|�0��$(�`�vvͦө�Sp���,Z��U��
;guWA���e�Q��t��[��!�.Q^���I<I"0/?A��o��j�yp���!��%S�f�XK�������I19;Vi!s�~}���D��x��&��th.�ՎO匂N_w��[��x�� �G8֡��㪩���A�w6�E@�e��������!���iKfw���]�vz�}p�Ov�f#@ a�Q`	��	8�������3[�Qe�5f�Z˔L'+��-�U�D�}'��,���b�Q��ϷY^A8�5��Y�u��UV`/�l���j�fG�1U�A�U����'oVd�`r