��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L��w.�g@]�4��V����ErsHX.;<D�6܀@k����(5sj��D���Gн�,푲�h�u�x_�S5Q��}^�!��L sUq� F���n����@������%PQ��q0���Ή�} �G����g��^i6����R�a�J-	>�F�6�%�:�8��v��f��zDVGPzUsc��Wַ��e�^ݝK�vV�n���]�b?uu�}Յ�+1���i׏ф�(tIs;l������I]fS�*�cgL��W�b�s��Z0~��W�������� ���A%�#���O*�gv��71�ٿ�%�QY���ٹ2���![��lq��BiKӏ� E����$�C��l�\����r��u�^}<�A/�� �9���Q�O9c���5�mM��NkB�]�1}c�)��n����'���G��N��f!H�<ba�8Zò� �v.,�c�� �1�|D^3T6-��wm�("��ܾϜ����(>��ſ�-��%�D��Jh�A�70`N�y3=UU�=f?�徭V�<̭�]K7�p�G���$�Z��\5�{
�1�)HO��H���������kd�Ou��V?� �W�@���NO��;�f�'�>�jJ>t6�����f�^Hh�#��\YX���Q���L��ф�D/�1��]m̥?���G�zܲM�N�>��z��6�%������R��5z�3!!���yu[EM$<�����zz�b:e�K�-�@Ӹi_U��?�[��ypN2[3=du�&�=+�}x/f̹	����k�L���)L;�%�U��F;|��w���� ��fȴ�W���N��g9�?�gw��u=��a�w�ο\����� ��`{�wZ+�떥�<�hW&��-28r�4��E�?i�#|�H�Q�t֑��(�R|S4N�����<�k��n%wʈ�&���r�7vu݄
���7�G���TW|�%V�TV��ƌ�Кp��%��&��gvZ��G��t_�����\D�w��B«G�TўQ����V��Q��۟i���rT�,Jy�����[�����`�I���X���!KnSm��܅�\{F�^ۋｬ�	�6���0ֿ�l���^l��Thf��c��`kf��d�

�ߦ�V([b���8��ڶ���P�&�^��(:�)�mf�g�gk�TZl��֧	�_�	��pj6�!�m0�~�5C��-���J���aXc�3~FmC�A�]q����ϧLF}���ݘ�(4�3��:���5�J���@}��`�tQ��Wul�xL�%+�������	߅�����p܆�#��eV;���Y+���B�,j���^��J�ngb�@8]~}~��R��@�d��P63�ՠ9���!m�76��;�P+0/�n泀'�+����ӂ�+^�H
jĬQtU���v^F��ۅ6E#5v}�2e�Lai'.e�I���J]))3���Sb,��+�!���Rd_�
�����~㑕;I-i�'�ś�=;�|�w6W}��tA��V'{o��s'�:L�F�Ř�>�C�6F�����\i'��T^P3�ʜ}��]6��{�ͪ[n������Ԟ�D��<e�"���D���|;ϰK̗�M�$���[�ʷ]���S��)**��,q��Ս/� �!����K�7Z�
���$�+ ��GQ�����N�8r����E�R����s���U�ςW�-�Fg��B�n�	Ѹ�I&��{�q��kgu���0B"ةߦ�{��3����D��!.^���&teDhb�/��i���qQ���ށ�9c�Y���k�Wmپ6X�RdK��ߺk�XiB