��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<����6��V�M��k�Q��e=N��G�7�/�'�!+�/�����c?�<��N��}Ŀ��̸����8���T����4UV��A��b�u��D�':��X��vo��\�L��K�׀�`g��"f��˸y2�m~Xe���,�r�:i���1����&�ɠ,� ��?��X]�w��>��� ��#Y���)����ϥ�J�[J�J�%Sf���U;�F3L6���e9Ync�E��5�Nm�:��D�]��z�/r+��)xyT~fsSZ
A�]bC��>!�����-�|�{~�~�\%"�7E�Ԭ0��挖�ZB��N���?'���!9�]��O�(���☫���:�h��&�/�~�� z�]��
鞊rv@��Q	+��nRI�P�W�Wsn��U��Y�J2�f���N���8�r����n�%�97{]�-qt���X���<�N;nT�rUn]�)ˏ���\���֔��������	.SP`��z_�@�}��nΝ�����q����.�fOIl���c���X���m)]�T@"{
�
.2˞�?��M�������f٧�U����	a�ԶON6�d%V�Epc1:#	����M��~�&��H���ᔉFV�@]��%'��2�;�����6��z{�q�W�3�:C/�W���+YOz�tU[�^��r��̢��u�������Dٷ��|�!���:a5�mp��C��>�Qrz�6j{R �3�u�+�9Sv+Y>��]9?uNm[�db�=���-'膑�-�,��Ц���v@�G�9�r��x��@JL��_����s��_�x�~��iP�~�N�J�+~;��ް@N����W��,N�0y�D@\ ��{����K�D��B訠!P��M����˥�$qH�1ѷ>����ݒ�J953�E�+�2÷([��� �O��Ae�9u�f�}�g�G[�GSAk��Љ*Y�F��%Tx�)�7��C��b��%�r�-�G|�$���X�2���咩�[��Sqʐ���u1�p�jK0>3��P �8��1Z2�o���V�l���[�yf��Z�3��s)ȉ��Q��8sg�V!Y{��Q��l�M;��aM�-�-���.8�������ǐ���v����UBM/��W|w���Q�z�}�.s��ge��� M���z���=�����3E�g�U�YB�W�C�����G_�{�~L���y�.Q��Ϳo����p�e�gI:p�9$�)ίP̅o2K������#�S��i��8��YM1�ED
�ap����A'�NB����{�I���<>b��"YԎ�r�I��:���=�Ԏ�b�j�M��~���퀔�P��)x��\���p�\6X�B���<mqшNR��>cL�^WS&(��$�c�k.�ôT�eI';��6��\i�~w�����+ǜ�UZɛvG�>7�z�����T���@M"��@v^|���Q��u��{�0���К��q�����K� _�\tAu	EE�T�����!���W��5/����˝͕��T�>���xu|�ۿ�Р::���隙�}T_��uΗ����d��4���'���)v͌�������/f��G�z�A�Y�|���+rc7EјX4t\�I��&�*�Kᇳ40���sK��i*��(�j�N�c�����As@���u �y�F�&hu�"��^��Yr���,�a¼�W�H���fpT���*�G�uX�_dO�5�lk�BkJH�[Cm�U}LT��(+�)�q�,#�F �,bKB�:��c�B�D�i�|