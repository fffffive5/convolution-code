��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<�*/��컆9�f)/�2��ڐR�w/���e>�SZ���kH��VI��0
mD��F���K;�p���I�4nfPK�>?�ϟ�WՇEIb?�(1�>A�sEZ���Ѡ���Z�����L�ym���>[��$������jS�$�l�F�8_�3P�����ۯ��p�R�a� ��")�ªYiJCW���|��R�<���EM֣�DV�ҵ�-׵� 6Q9=n���6�7�sP��{�R�=�9���tuk{Y�p��n⸰�+��M���y鏧�W��܇8� �Pw���_x r3ۻ8�$�c��=�|��\��$~��ؤ��'bu���@��ڥ�FP��]����ȪuT����1�u@4"�V\,bn�+����\&?G�}��v��<ݧ��[�}C+����.h���Í;�D)���!��#�Yz0�OY�;-�Fg�)���Job���لus'��z�SÕn�z&o@6��+�!Zd"ij�����6
�����(��\/��h?�GH���|�����"��k�&N��z��em)l���o��y׿�zՏ�(�}"z�I=��߹}͂��4c�Ne�,Cu6��ݻm�]q�U:<�_d����w��J5�в�V���ȏ>@�i@!@����V�B�4�͢U>CU�
��޽��,s�?�+#�MpQkO�O��쾤�q]��Kg��@5h��*z���Y4o���cҮ�%Z�<�G=���$;� >��)ɯ3�P�@��hQP��8�#f?�����]�=LfѬv4�P�ӝ�~	����=ˠ(���� ������KlڐϿS�6�'u6ȑ��7`Umb��������$E����aY�o\huo�A�� T���,�,�G\����v�_4�"K���{*uUm��U��ȠZ#BV�eۨd�M�M���un�����-�C���5���uW��v���>b��Lj���|����z�u0��N�M��pd1J�+?Ա������1��
� �=<�^� ���`�+	�8$� �Nz>{��&w���Rp��}5&�lUKd����Lͅ�"Ogҋ���9�`ۀ@��1'���S�����wp����`L~�H§:(tѳz��&c�@����Z?��*�?�R�7'�@W�$�d
S���o��.�H����7����aJ��*�B�>��R�&rB�0���~�ْ���#`�M�z�Pʞev5��x���LA��}�	�`����f�V���^�J������ʊ���N���˭���>��B*\ ���ݟ �3���N����T�j�����`�s�h	$e>򞲓'[j����~J��1ޡ���F���TB�����^�t [H*�B����6�&- �yr|�(ȵ��@�Z�^�u��nD�y����gh5��-��r�9H�� �҉|u�ku}�Cn�&q�<5�&�s����/��#k�1S�jb6	d��adv����@�	W�$��+<F�R	xN��Kωr��H���"Tz�=�ۛ�Fut���&6{w3sFO*�/=�j��^��I����u���(O\������I�G0M�^���§�ѺAs�r�X-)CN#�>&i�Q��ҠWp������tv4z���ƫc����er��|u�&ٹ�<��H��,k��Җ
���-H|�>Á�9�?�_4L�}���Y�R"�u}� (���)Q6ڴ�0qk>ɺW�.{�ñWc��%��V�X�|��k*m10��}E�s���A�S)��[\/T�K���!��	���k�u�Q�<7��{
�3q���ڄW�%�T4�sPw�t�Yt=U�P#\�mQ΂�TaVK�=1+���-�e�k;�j`��ܞUi�o���n�{_��Z�	V�i\OI���m�\�5[eĥ@W}�ɓl���(�v
���J�匿3n�̨0��L�����5��N��ezip<�-l��K��o����c��T�t�"�ߨ���>N�*�nfõ�͔���fjq�m����hZ�ˮ<7�:b>���ءלc��F�SH�Le<�h@	K�7�s��i@��J���~~OA�'�,���f�7c
Ą0��h6r2�]y���&+�L��o�&��
A�9���t��*8x�f>V�nV+�VDKp�{��f0�� 2ҝC��P�1��"�<�!V����6̀[�ŉ��^�A(~�1�cQ��J�tҡ�BƔ�Ɋ` �0�hz���$��X�Χ.#��w�8���r���i��hl�t\�u[_�)�Z��,�PzqL�VLx�� ���K��ȹ=���G$U��
3��8س�g1��zϑM��$�҂k/%Q�O��K{�&�"�6�l�5˴~�	��f���Yj&i_,��������'ԛf��@�6X�5�Y�W��S�$>�]ZA꣦�]?�RT�4��/��j��S����Zx0��r~9� �XҿIj�N�e��T�#$?��*8QU�vд�� �o���//8E_N붽IxG9OK���e�����RA��%RKF��4��/����Q��C,#��q�����l�Qf|�Lˎ�����jƒ<#�� �u7�M0t8�LW$:�S}�����B�\��>^/�l��	|2G7(���\�Y���D%��F"w*�z�WmP��@j��9f�^Jg!�K��ˍ1[���k�R_*Ԓ�.L�z�Qh�`��|�R���X,N��k��Nl�`;F��g���B�H	-�G���鰹m�Ɍ�m˭�ь�`WfqU��ǅ&��K�*aC�:$]�,�?�rx�OQٳ�9��w�`��>���`��c�~�jܬXf�	܌T�t��6đ85�W)��ޢO���>P��QT�������R�Y�V]�#L��	o<��8�)2��j/��T�0$4��N��o�>7ɷ�ڊ����"}}����_~�5?�{Y���}��O�e��I��]6b9얼ŶP	�Jj��o�a�FcS��w��s�]uck'�
ʱ�m9ਆTL�m���$ʒ{�U� `A�-�J4�OgdkC���y8q{��H+K}6��Эf�c�������j��UGp-����W)v{�=�-j�������,��*����[��<��IG��yu�(J+?�&�o^��j�]��=�1�1=�]���ϓ�h��m@�DL��ؓ_�:��qx6A��a�+Dڋ�}Q�]4�ݟ�ph��v��V�V�{�0�F}�yZ�c�U�ĩf���-�Y��8���ÛG�<}"lg9wnʩ�{�
k�=�x�T��f�)xS�X�`�r��#�w�����H+�uB�E�}�q���* ��U � C�G�\����X�$�q|�)��y�@�§�z'�-�j]5=Ƌ*Yףwmg�n"�G��yF����t���K�Ȅ���jp·����,n�\[�q��,�1������r=l����y�x�f��OKn*IR:��]Ƒ;:�����^�5v�L���L�ϒ�h�sa���/"�O/�>��6A�Lw1{λӜ�T�~w�]i�eD�ί��Θ�4eٛx ��r��f����Ņ��I�A%�ɪt�络�|����6�D��<��x�"V�:`��1�!n���
�	��ɒ`�0��!��9�n��{m�k��6Ԗ�]�@͗w����`8�h�ֶ	��R�>�]��p�&ȭy.S�f�L��ۥ
I�Ԅ�b��r-<D����dO"�+�f� m��XQ�#�.����B�B�媑Gh*�sY�%W�z����o��0]��i:�ۅ�&�4�k�]I8�A��^�����rg����,�7Δ̗��4?tJ	��]}��ҩҢ;��"��ɚK&��ΈAN�޿�^|����rz��ZX!��運��<jO 1쪲���WHJ:��4�����3�Hա�Y��F��o\�!�U�����tc�a4$����(�P�p���G��&��r��ݱ�h�~�x�Km�r�c�9򦙤f�/Aw�CSB�3Ƒ�493����Is�;�Ik�Y�P�;��j;�'CMVȆ���O��[�<��73F
:��LS �����a͢{|�C Ip���2�A&�&��O��*�U�2���������9�/^Z}����q����p�1�ONm9���y����q��&�b&�FW��u��c!F?������%�iQ�03���c���W~���;[�?�~�,�2��(+�q`6�T`��r؟%��Vk�>Q��3s�l��:0�CyTgZ���F}E(%>%t�`�[��U��_�3�X �����7�� j�����J&Bs�����8��]Ú��$����rTcE�%��`$~��1ܐV�1�GQ3Һh�<"��؄��.t��B!v�>=av��������:�eP��&='F�+�v��k	�R��A��c����=)C7��5 ��o.ʻM�
G����������j>�5���lnr�l����P�d/�x��Zx=i��˧u�ݬ��2ճQ@7���*�DPq$Du��J1g�X���7�\�^VqL��U�l��1D�"O&�ׂ���'����Yz�=�̈́�$������YK�rjb���ڈ����ϯu��$1�%�	1��!h�v��@�JYY���.G�Z�y�����gl��^^������FS�k���]���p�[�2I����´�1�Y���G�iK�iQ\ �E��>(����
��[���7uf�I�D�rC$򘠗}!'��[�oq��+I-,�C�7�wBL8�׼���Y~�>����FN3���0zr��F�3��*��_��40}_ⷝ���ݗ��l�$F��N%Wc4k4W�jlv�`��p�L?�� ���?�m�\�C��Vj���r����-L�lb��p�WH�9��d*���׾�F�bt�A��m�'(-I����m~b�|�d����N
<��o�����6E<�E�Xk4Y�I���{��=�X��	!l����w�}p�W�:��r	P�:)�]|��օ���}-V���G��
f;��:��:I�~�d쭆rv���ڙۛOwD���t�d�C_�����/��N�a��>,OM�cSa�B������?$���!a�L#��PVI�����`�p��)�(�7W޻��]�"7�Ae����[�R��^��2�y�|�3��J����!�Ӵ����'��C�.�ƛ��ۤ�ǣ�[���1�L]��y��S�Z�4���C���]�&-8V�nT�6<wF��4F���s[A/�T�@miNǟ�7������L�%U������B�T�����{Z�%&Y
��X[�=��ngϤ��W�jyk;����0�9�^HUm�'����DN�չ����J=w�g�5,��,?ɌU��8��h�����G�	u�0�b_J24�<o�G�k�W�Pdl�v2�6{OӶ�����*I��T����M�1w��8�� Ŀ3ݿ0n$�_�*F�ێ���W�Bj�������������$zq+v%+�j����fFbV��)�,"
@� ����d�#���Jd;��L_2����2��%�A�˥g��;�f2����|�L'`�S��vpJ�y���$��]�'��h�#yF[��;_�`V������9��-��*�W(��E������j�G,��1}�SwQy�^,N@u����O(����f9��([p��͈+�}ӕ1���z�|��h=�����\�]��h))3XB�/���w�p6�m��GTH���S�<��j�{I���l��a� �4����*�̇�)�9<\guÜ�`~�qECn.��j
������_pܣy�e���}*I
�B�y'�zr�!���ה�GGzE��?�n�.��%VXw� ^�ȈR9�m���+�������)w�Q�x6�o��E&`a���'WT�*%�Q�X�����0�}m��&(.d�_E��E�M��v����z-�[A"r%�|_�е�0/t�*��q˫�pv*v�:�fNlųJ�qw�V7�D��d�:��=��7�Xi*	�v�X�XU��
���YI�S��m�;����x��OV��kq�J��@�c��3�=��ĺ�R;����/Mݤק?`�N��2�����:ô�ѝ��^�sRaXC�0�Qn�le�L�~S	�v��^��`P�>Q@a���R-�In`/|� 16�nR�ː��Q��,Jg�	?{���8���^�4���Rj�6h����l%��Lч����N��N��O�����	�!O��?�zj�����<��u\�i�4�<#�e���CP�+O�v�p5��<K�gY�?�5@�b� �gC�D:Ƚ'?�߀��ӝ_-��x���Y����+E'����F�w�BbO]���\��F2u���)ulLn@&pe�h�qhB�6R��[^)WV���j��΋�C�0J8�k/�H�oj���z�-/���Y�ج�̼3P�,MZ�n���_$z�={��͊b�`����1@��� ��	[{Z�݇`�cX��$��ǿ2Z�wQ���+���d����|	� j�:�]��Oі���_Ԍ�������B�b亯���%�����ȹ0r���N�xh���u-n;�)}�B��F'GΞ�xIx����;�^E3���	o�וG�$&s�~�#�B_�*k��j�T��D^��w�z]^7~�m��'�?��V?���n�O��f�Z����5K��I��T��51�z�����6�Ƚ�'TIґ��B7U2��~������EV��{�kF�;���@���ΐ��ә@�g�%�i~�a���DJ�ϖ1�� ��5�P��bPMDN����Vr��%.
���m�;��U~-�yK���፩2>�}��q�IK��,VC��I�c�|!f�~M�"w���tge�fK�0��O�ғ}��8靿�X��&���R�/��&�z�O� ���Vg�݄����Pvi��K ��Ywxb$iۦ�����ފ��{\���_��A�-�<6=��[�Ѝ\�k?f0�H
�J��V��_Oﾏ��$$6�ε��-��▝wc��>mpx�G	�Q�Ũ>i��"�wy����Yہ;.�ՀɆ�z���i'F��۾�/&lPD"��Z��GR�)�K�l�l��:%���M�mC���hڮ�T#��l�2Ȇ���u>�Eʮ9r�E�6a �r܃�������t���m�E9j�euByJ��9Y�����v�̸�SS_v\��!������XV�
TX��RI�]�\:\@�"�7���+y�<���%����b�q��������9���������hbϩ�V�s����WF��3���yA�ސ���0��IY�'f7.ΓE�U�t&��ԘY�*���j��k���s
��@S1,H��}w�/˴��[Ns�S��lU�%�����m�S�!a	��=������A��S@D�Ά��m�],nqi���S켋@�K ��L�hB�0�A�����H��j���!�e�����k�����}#v��Z�3�|6G�0'V�ʖx�G^P��}Ƙ�e@�e����E/e���s�LD(x}ͨ�a-��*ũe4�w ����8R��Cًn�ȕ��?��G�����'���"�� ����M�(?�0�׍Z�I7�ԊXt���~�%ZLߧ�EW4��6G�'��?+����D�`1-��wEf��X���,�N����Vɤ�T��i1���.���-;]�5MO�gD籹���R���IVRC]5�r�w�K9���浂`%Yra�j��fL�}	QI	~��(I���	�m��6<��ݸ2��^1�ؐJ�$���v�?z��y�v�e��G����}����H���֭��\c�q�J1tχ�4�W��wď"���5���n���6���dc�_��������%�}֒h�=��)ўS�f:s�/�a�O�3��[SZfuި@���`s~o���d(5
LzX���i�m��!�ΤJo�����ʉ&\�VN����	�'�Ť*�����82��GpNU��(~H�(��9�蹷�� �4w�8�k��Lu߂T��v��:*�	��!,��K�����`o\9W��g(�c��ш��.�p�uQ�m��tO ��b��I�+�����+It�:�T��b����6�g�2�r�)��_PO��r&�O�[.S�9��t�I���ct˺x��7l��ʿ"�VFᦧ�Y���>�G��z�$�����s�֜iZX���f Vo�s����bp6��
�Jm.-����A�ޡ5�h��H�u��-�l�(�ϦL!�_I��'�NI�S0��� �K�3\
]�nT��FϿ��U���R(��SH���TE�z��@rOA�n$k���=��2�K������A-r�l������2P�J��b(oڭPYy���GYQx�Z-�: �͙�?� ;�6�7���)�����v��-�o6��(X��⁦�k$���VF>�`U����6cOgn�H���F�B7�^(����h��"��J_02���LG�
I�^���R�.>�{I6 #6����S��5�T�pIȶ�+��	���R{��t��b�p����ks(�[����tT|�/����T1w�Γ̀o.�}�����]�ܢ����Ή��s^��)G��{����$�I�J:4��CI�X�R��֗���W�����ڄ޴�c�FVȈη���_��y^��G�@޳:,�7�2�	�p\% 9�,x�C�������#�� ^ۙ���Td��R���E�]��,G�2�%�^�[�FE���q�=���ߴ��&mf�����2�ؾ�߽��t��)'*8TD�/eU��6�n����ó�#�E�=߾����Ik
*��:r���a�T�6 ��4�����Io�G��g�PFc�,�<["Ȣ�mRL��LGY
."���4�β~��hn�q`��m����}Ϧ��U1�\�1q�PI/��s�T�c�y�fQ�Kd�C�U|�N�;�@��t��I�Z���n�!�[wR^��X��ߕ
L�D�w��������<k�}���˴nfy`>�ؚ���ㄌՂK�[�`ۻ���,�i����nfm�Jq#������3fj�b$����3�W��� �HhH��}��	�W�Y�ZDi�2���vۂ��Q�΅��:�[#بr�Z.�0w�n����;�Q5���ĸ�a�X���Ea��nEW�RN�W[�U~����#��tkR'��'�.Eq����8{��U��˼U�@�MxIeٖ7Wٶ�MKJ���z�U�!.�{m�A����E�Q�`�ϔ�7�濈ԯE��O��Q���c�}8����	+$�W�/�$<��Zl/ŗZ��9
�P��گ#X���=�ns�JG.����rs+ssT��H�2��Qg(J�2s�x	e�	V���&eY�,�{�X�K�>��Jo��j'���'��Hr�<U��u�W��������d;���^ۄ˙��9e�A
0c-ŋV��A$c2����GB�RR�"7޸H��(k[�\ه�s`�cQ�Aj�J4���%���
&�F�G�c�?0H����ʈ�2>�^DXN~�-e�v%1D`��IL�aU��*�.#�H��%����Qc�xY��Q x+ ��H��X#`�s{j�kx�dS=��R��&��0�>������"��o1(/R`��t��A�n�v��YR��<=���O�O�t[�e����m|��1ȳR�;�_���7v��Q�|6Y�Q�l�9p�ng�K��p�e�n&�q} �����Uwf@1�R=7u#����5b�ĔaM�&�;8�0��;K�q�)㽞�������<�l�޼��n$�t7������k����=8S����1�p웍�������}��@D�Zx�Mr���A�Z(�٧H���d�����C
Odz*�`Mǂ��K���<;e�a��6�i�h�B�[H
���֞��f[)� �vc���+a���A��n��#t�HBg�=:1wB�����å��⥁v��_{AY:�T�(�'��P�A���D��?����@���IX@�]��8hQ�+��X�	9/
d|�0�N_�f��x�!�;�|�qv_HGj��j(�*��7/{a��U,���o���?������d���ia����Ur��D�J�b#d<�Y*%n��D�Ŀ)LD笒�k~ xE�׾U\��0/�:l��3g�Ώ>	��[>�a	S���m�hC�/��!����C�V��O�����I�?��BYh�H�[��lԫ*f��[My��h�Gs��{���8���v�<���D��h{��Xhr�@��J�RNe K�n���l�8�3�-XQ�nc��ׁR���`����e��Y��-�GF��)�6q�a͡��K�S���'x�H\S^�y�r݁����RB����zǗZdt���ԺP��v�;fʐ����:^(�Iٴm���&:.��j���pF��]��d��[�r�̮���oj�.�תS�	��G�S�蜐-YD��.�s�ٖ@jD�7[��.�%K.W�o�&M�r�n��Py�*L��NI���Ἂ���8Q�gY%�|��׳�u�o�``���6�O�v����5*N�d |:��[Go=G8|ED�6�� ���?P�j��e��>qW�[�W��E���R'Dn�ZJ=�a�g����gT��bw�x�H�	�`�������.�EDfݥ|妚�+G���q�@�V�PCB�;�%`(2l7��������&�-��-d{�ps�ħ.�ʈ	���1e׽V��H�d8�M�D�m 9�m��gن�&���L���5������Q���H�W�&�姢q-��J�D��-Y)S3��d&NBR}���>g&ka����J�������Fn� H��"�ϨӨ'ў�G%. �VXh��Ϝd���|�^��y+Kh<����bU��X��5�@}�9����VP ���pըTP�8���#j��yZ�HfL9Λ|;����|�/�8��R>S\	D�Ԭ�֖4�K&�q��C� �\AIB�8�
�&�TܼVvy�Q�b����E��W�M�".)LI��M�c���:�zˑ��R�x�����91� oF�tE
��'p]����Ho��V	[����1FA�l/f-ϹB�B�"�� ���������DR$N� �3!�t�?�g�5��i�Kir�j=����X�Ϩ,������^���bޫ��j���p��Lj^�����s�lRw:��˫F��x;�x$���2yh/!�n�9�L�b�a��Z��<_���H�)np>��0�K%%^�ˢa�)�:���xN�PcK�@������F�%�^����OC��ؔ�;,��Q�\g�-����
�`����~���iS��-xRD�ͬ85�R+���~�Ëc?�,���lg`��Zs�Lv`����W�wj)l�ӱ`iplg�J�$(��W�����_�,T���6��u����6R	й�@V���G���sg�Dq�}���}��9c��.*«��BO'Ԕ�ǚ���
v,6�=󸹾���Б�r40�����IQ?~V&�(�[��_�$	���3*��]�	WBj�*����D��ҮaU�qYm/ �0rh5#���1�Z��s�,�Fcf(��
�V�����$�So���]�&[��G�J;D2�]٢�,1o'�a?��͂�A��q� m١tƿ�Q�������/��q7ϑ�RA㟝�{��G�Y��2|��_|h0A��,ʞ���t�0���/�(}�d�����nk�J_��7Էl{Ev��Po�е���&C�ǧ���7���Y�I�T��R�?q+Y`�͐���,v�Xx8�5D�u�n�I]��甕�刲Ʒ���~���b�7Q}��[����F��uÛI�Ь�a��pf��;�c�Tz [j��3�