��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L����ʩv�*z��(zH�IK��'�����g��N8�Y��!��*	S��=����!�@���� ��׺�5�/���d�iЁ�qb�Y�b�~n� L?ګ���T}`�p�::�D+)�\���V٠���^��O@Z��y?�SՌ=0))�גE��2��3H�$�=��]щ���b
�����T�5(��5�@���'��Eø���/�%��&�B���F�om��X�(ۨ��^�M��S1�,�״�O̨�z�;V����w?�XHɇAj�[��9����<��h��0���+����Rs�Q��- ��2� ��0�XX�B*+Iw���$�������;W�]��U�"�{+����Wx�)��
�5���TS�����R�KC�7���Y�H�`0�>�!���U�Z���l�P�������sh�ؐ���ي7�ާ��N�0Y?��c/�L�H�%�ҥ�Fw�?�V����^vBK!�>���dp<�1C����)�����kg<�]���8�&��n�w��i�H$(l!aZApɬ�Y����#:���` ��[,w)J�%�SarǮ���D�͙+x�D�re�~�)��^ݲ��Xϩ&U6L��x�t@��=���}3m0�I3��c1mZ��XGc�pf�4�$G�l	K�V"�g�^t5O��cW�ie�b����.�gv�XA/��?��b%�=�8}|o뱙�AWt��6���j���O;Xlٖbw��1U��X��F�� CT>��>��e��1�q�2��fok55��OO|�t��k���xZ�Z��{��A\)�k��g4��8�L�eTu�^R���d���@���������=�4��A���U��N�`��g�j��dN�۱i�ؙb�׾l�L���q�In͖��3����I 4�-&j9%�^��P����u�uXH�&�����l9�>4�z:�-�,8���������ۯ�r�JA���*�w'j���zNr;�1��t�p#Ȑw�l9D;�iD�@e����1���3J�����j���R䣫���c��r���[=����yt�/TR������b�|�����������g�lwZ�?�����y+��T��'�5'>������@J�������=���SZ�R7�X���ℓm\�Nq�]�/��eA�!<�O����JM</U�t�F�c/�}cu�6��'!GD�Fy˒L�Э �c	+8�8�|c`D�m�4@��yo����i��$.&q�����<z!�߅���F�{�ܬ_qԶI��Ԥ2�(�E&C\��hĮ74�ԋv4(2�F(�-�6h���Z��+4B^]�%����NbYޛ��]Y�W�C�"W���Ha��  Iޒ]����>N[���`���(9n��15�^0.�n[9�̶4E󓡠?�3�ޓEK�:�J4�ڮ�V��5�����U��0�ov;�-T��Ւn�R��Wa@��ोDA�v4/�X�?	BĈLϮ:贁o'@�g��j��H9�"&Zrtߖx}��=���6��'� �%��ݖ3�� cɳY�`�9q#��W��,�%�'��0Ա	;S��}t�<�U����|���{���na Q�,�~�2�b	t���VM�V1,��'���Vk��$�O�ܒH����]&�B��ōa3�*����ү��^����#±[�`�$��|�>M��Z�E���qX17`}��4R#᳑��ŷ�]+�s���I>ϗ׹ K�޲��7V����me�E��:!�чI_2\��E�\r�H\���g! S�1}�1��!"=��,]I:�:�J$d�6�ޱ�;Ww��& )>���^Ҥh��&
�9��ꔅ���=|�P��/J鵬"~ ��r�h�MQU~�s��_9 ��	���Ood���є7)J�:/���D���XS�7}ӊ"M���.��2��\i��ا�C��F�w5+���߉�^��/���i%�ފ�[���xq���F���*0��3�[/�d��L���ݥ)A�c�*��y�:z��r~�=�2�}c�uh��h�G�'��$hc�v�Vd%v�C�`�]p�=a��E�4��b��,?��q����3�C��E���Z�]����7e>�_y���§���Leo6,�N�*p0 M<ϹE��"���xϡ����	����/��G��C�7z��N��6���&�y�#'��VqU��nE�h �+i��J%ꞏ�|<�Ȑ ��@M#�m��7��+G.�+P3ڱ���Z�()?D.�E��y�c��@>���'�����B���tF��e^H�ݐ���_p	����kj)x`�t�l,ˏ�G�r�J���
�Nb�a��\r
�y#DA��NG�K[3m�iaw�l��k{$,�݌0Y���HT��z�aXw����ۑ��@��oxY�h��b��>&8W-������$��>o�K[2��bv0��HF�zm��=2�ȁ�&:3�����?��ݐ#u�Lwj�j?kȁ./��h6��sqa���w>�s7�
�YU�[ m?���A^�k�wa~�	����[H��t�-n���vbLG�k{!�G�.�&��`T
BAfr�����3N9��l���:|J-�?D�k���_�lm��z��A�Hछ�ɿu&H�����\g���P��?G\�g}`g���kxv�[�F�M	�%���:���\Gx��ܟ�x=���MZa1����9��}���R�}��! 
��p�s�J��ej�/�{u[q#?�M�7��D�7��g����7��&\�xǲ
�쏹�Z%kS��l�N�)����gAUаb�5�R
�ĹXz#�h�8�ܚ�2f��e�$%�-)�����(�Y��Tsy"^�
��hO�fv���?יP�t�T�E���d���&�\N�H�Peޱ,Nk�M�Z{xv�oI>q�s�}>��C-�Z%����q,F��s�:N�"�5=nsj�f����j$��*��쒬p��4`�k�^������$4 -�
L�-�΄���d :�h��\,�o��'B�y�$�U:w�O��_ŵ8��F�!_a���`?|lYhY�����}����K��0Rz�[�S�F��-w���+���W�Dv]E���r�t�j�a�2�R#���029���Lw����,���$R.wWٹ&����{A���l�a���_+��)�)��(�x�D9d��^eyv�ڛ:��AE��X����&{��=��ۇZ9"�����k�B�:�
0 ����H��v���?)��t�J��M�ǻY�����i��UVL�QѤ��	V�^�G�ݔw(�0�q5���k�nv"���Lb������vd��.�ɭs��u�O����x;��{O�?�e��K�i軀�:pح��q�2�U���#q�&5Lً<�OL-�����
q�EcɿҨ�u��/�K����\��n��l;K���������$t!Y�u�E�ħan�ɷTY/k9�+�*C�L�{�?9�=��er�`L3�=TSJ����t�� ����8]�L%1���{8@4�i�e��f˳�Wd��	����"�ѷ�:�� ]�	��\^��Ȱ����"�J���DdLe�9jl��u3=��%1�@�(r�n�3O� �.Ь����ʧw����j���b��&.�\9��hR+Q4�D?C�.���NWT�wxJ`�LQ"�&��$�S��8��:t���߷
t���mF.H')9Y�)�X�{��(�aN�|И�9��Ua�GG�"���9���Fh[
mO�������WCE�F )\FL�j�O�U*����5q��Eb�[c<�I��5]����⻪���UAX�G�,w*9Š��M5b:���O�i1�;��x�%T_�@=�YMb������թI#mjm�3j��:K�+hH&鏊�PC��N d�I;�ˎ�����;�0Y[�D���F�&�d������m�ʮ6���ne�`�'�E��k�Cy��|Z/"{��d�^����8�A���q����e冄�f��+���'�=�/n/Ȗu?z�"�'��#	C��'w/�#�D[�J��}6\h��2$�h��
O��9�q�N|��K�0D�7:?���1�aa�?͉\,�q�䠈Y�#I�&7�ǚ ���F��p�C��+)�z��H�=��ܣo�A�V�3�>��^D0g�26��xp��V�ς
�;�����v��ԨK4&D>�:[����dJ+�խ��RT`�`"�Q��Qsnf(�(�f���������Uַ`�|�?�-y薐����_>ǔ-h�f����Ԉ�=c,�ܳtx��>�몇ϧ̽���m��L���aQݕ��j�~�ԋ�%X��rW�$�{ޯ�z҄ҪZ|�b�Ye���رre(�W��o����U`PmK.<�'�B=X�Zu	����@*��ǚ�x���p� �����oi���l���˒=��5��|J���s��� ���q�SQ	c^[���u+l��W=���`�r���50�~D���Er�:ߑM�ʗO�g��̌��\��7߮pXY���:i���Xu�~" E5a:'�����p�~�y����
��t�1kE�`�1���Q�Љ��p��Fӈg|�T�Y���`ɾ���RИ�cZ$��s����q���뉞M�A� ����d�^7��Z�������u��t&(�s��'s��j�;��q���dO��
����	yfd:V~���e!��0iī�v������[i�*��p쟘O�t���d�Ϭs�x6�E&6���+��D;�B��ZE0:I9�X��z�Kf �e�Jm�e���Ol�2�"�i-�`����%�0nU)�a�[g�9�ʤ�B�/uZ�2u2����)ܻv�"���(=K03�$?Je^ �Q��6�B�*��G�W��)���+�F���y,����O7-|#Ķ�W��`�	#v�%+	��1�~�@�-�cMw��܉���m\�UR���o�s�3q)P>�ti��Ulu̉�����\�5����U�����y����º�.g&b�MeD9�[B��%*!�\���xLF�K�=���'U����o�*ч�[#'p\h|n)J�������˚=?-��!�J����[�(C馉��02J��T�J��Q�����0D���/��?oK��7�&����$�_�2��rQp�|�Vg�� �ŽFW��s?��l�Z�����1�ՃE��b�B۸.n鬦�̌��{zh<H�1�C�;�l��ti�E�����S����Z��˘��e�I�üf���6?2ۦ��e|��'փ=��E��u�W���?]�yE���y�Y�I�J�»6hk��ȶ2���j��XS�+^̫d
Do��Ԋ$x�f���4,�D_�;F���5z�m~�a�Vx/�	?��(ݡ��b޾��B�r�+���î�g�S�O�#�>m�\�;'&4��i�b�������B���6�rC���@F
FO���-�p.+?Iٗ��V�U��)�I��q�V!�\��y6���{�8e�����8I���ͤ|NV5k��Ѐ"U����s�>��'U��Ƞj����Tj& � �4��?fm��n�
�u�#��v�;��1�q�j��{a���Lx�DbR�
E��K_�4ګ���o����cׯ_l�cƑ{a�0�R�\"@1,�A(�[�]�e�������_�(�D�A���_)�]娖chk
hVW���4e�k�wL�%��%�L�=�vI-p����ɢ��`$�BC��w}������:��j��%o�>8�����6�����#V�ƀw:<��z}�e>�	�e�o �j�Q��$�d'���s/*t���^���p��+��~�[�7Ri���}λ�𕸓�bf����q��}%���v�Q!S�HA����=���JA�T#hU=<��9�O[=bCs�6!���BNn��Ɖקj	k�Զ|;��5��$?'�W�j�{�4����(ka�Co��;�e� 5bݥv���;�O�����D����;\>��CO��l�"�xw YdQ�,3c6��-���r�5��"daY��e-�8�a��5>f\Ip}�/��:ukmH�C�����U��'-�zWG\ �ۥI�^�nf�SɬXm�Bb�c8%Et7�x��U������2r�:t�=�ۉ!�r�ă�֍�� <�m@e��1o�q���A.�04�[,�4�Q ��h�}�,\s��vL�(��.*u�-�TM俐���lK��#��
��;�k��=�~$ �^>����!�)G�+�Ĥ6[�c��ˋ�SAseb�*;���fD1�,_�?R�+���P[?uB]0M��k����c����&�L�6�����Gy�*��$1�%�z8�ʵ��R�:���	~`��n�@�bb����A�D����8hcy���n6���`RI�]!�7��3͹��h;�뻘���s= ��}5p!��"��}]j�������m)�s��b��(���'���E�5�7e]cE3��/7NTtC���.�\A���s���xH����C"��@]{���?x9� ���@e��p^y>���U�n��3O>h�DE�Y��!S��?J��!A�y�7�C�
���F���t��Qoo��D�t/�_���qk|�-ؖ@�� ���׀I�~-!/�"��r�]z>+Z�w�3�[>�s�2�9!�%v��Y�
���{>7E$�,>Xޗ��F��]�ϋ��W���D]�3�F�͐�ô��F��4i:#��ȆG�ޛ�a��~e�ϧ����e�FGe�c�I��;ߕ\�@N9 �%�G��	�.Z�}���kA8�#<R�Z���'��.�C]/�٭*Y�͝����Ԅ���w� ��U�̖��'���l!]��v����F�!g0�b??
�U�Ȣ:fZ�����8:�f���+�<�����fj�sI�jY[z����9��s�T��q/}�K�z�%=H�����ҍ~?�V��D��U�l����yM�v�& �����nA�4\=��4�Hg�<	���3�N!��;�ؕ��u)�|����=
��!H�uCx:3D�����gs U��|i���/�I_��FV���e�=�5�3��%S��m�m#Y�b�����=��.�W_<�;��ֺ߬3����|���r/�41'��su��4��M^d{d�XҠ��E�5�:��q1�w��O[Q-��Б!�j��?&��,`n�њ��7bJ��ŋ��cA��K�%�`�n����@UA5��b8��a>�e;��9�x�.���p=��p���n?�h����,���!�٧5��/�l��[���4"��6!!�I�C~�C��g����ݱg�>�j��L�(l�������d��f�O�����t?�,�sl�j�ʏA�톔ŧ<B�eXv�ڊ�X%깪f/,��OP(�,�@�_�$��ƚ�"�+�=h�ha���R/_�әl��4�Ah�����l����gC����O]�]e>u��0��.��������b��+Վ\<Ut�+����~a��훏/��=��5 �	�WT����9��Y;aq7��ɥ��D3E����1x�y�"�PvI4������]�h��_��@o��ɹ�}Ȓ�>!f�#�
����=\���:�F25	џ�]�g�'"GA�m�4\�^�B�z�\X��<b���lQ�w`��������5Z�6h��d���oG=xGTL�J�,�+�?��S����(`qh�|��ס�k7��D�+)NB������(�"cM~�^�oӭ+�
����po�/�$��Q�3*�3�8[C	�:k���7:�0������+��7��z�<�&�Y����w�6��zg������B#��[�L1l��cg0����V.V�o�_���. ��Gr����i��kU��h��5�cC�cJ>(��W����q!ϼ���� ƶ��ll,}jR-�=a4��,��yG쪐Q��`�چ�ʬݥ�y7	��C�p�8O�.K�I���Ү��B;�.�*���Ҡ���f�s�v*��A�5�h�:��v>�*������.�?EB�������E�S�q�ac��g��vD��y[M� �Іe"�VRR��W�%��`������%h�~�l��bQ�CݹzYw&V"����G)%�܏��T����0� K�PW�f�T�=��@io�;���qC�.���p�'��ǵ�g1l'���� -�����8�1~�+,��gҷ�Q��<����DW[�\z��wxaM���#����9��T��b�'oh����cn*=&;/d�Xb�#�G
k�jby��l3���
��)e3�J�(��#�A�Y5�JO����k�����AL%�djU_ve�;ﻖ���7���K���P�|��G��.�2k3��F���IΘck�U��%��m��xn�C��xd���k�] �c�|I�kTJ=^���넛}T���A���7k�*�髀2f��S�����E������W�󠇭�g76�a	eۙL�o	_)8�a(
��|t�$Gv޹+�⺓�d{���_���������������f�},�?�i/�I�	�ھ�W�@fѥcO\���&T��b��J��y��r�?��(^����#�.M�d�R}�Ƅ%&*�����+��rb��~N� �thYC����;C��:͘�M2�Tt�c�x�ui��!,?�fc�l֯]��2j�g&�1�2���D���i��a�ͮ�ƽ}���-�拳;�i$�卉$5M����}�\��#\�V��v	�T��B;��t�DR���%?5 _3���k�Ȝ����8�j	����E�U;�1C����Ɨ ����yM��dV� +��T�Ӛ}�6+�c�p���ؗ�^W�_��Oed�N��"�@�>
�Hٰ���=X� ����"绍#�͔W0Ȝ</��`
;���"��Ǎ�Tzzރű�;���X���t	�:���ڣ��^Գ��M�6$�~����	+�{��r�L��g���$���.�E�T���B��J��5�x�
ib������������H�I�����~���H��C�MO���~���O�w���&u�>����m��,��WҖ���o1������!C��w���NPD䶠��۟ 1��A�m�� ��6��N_��bC )���'��4��&��꘏�l�T�õ�Ӳi��|����L���Q�@��6n�����`�,��~���	�[������ԟ�y��y��A����w�W��Q�?^ȡ��N�8�Y��d�-�뮆|�d�/hbr��`m�m�w1��CH�h�qz+E�WKI�'�,}�Dp�4gn��7���;��;+����u~`(F~ԯ|��M�m���]��?;�����Sq������z��ھ#�V�^y��MÁ���Ke镄S�5�v����/)�Gي����$�R��8D3#8�uЀc*�����N�2�{��u-7���np��Ѷ���a	�����.�:��ūD������{���y�B�&��/mR�Kgp.�?��H9!K �@M�[KQ�-��k�;��G�۝��y,���	:�8�,Yu8�����P!ֺ���͉��X����]N�un��]��}X���'(!Y8�u�:����w���n��L�W��)\z�;�^PD�o���P^*"Q}^c>���_ܶ��Z'@]!�F��U�7D�X��N��Y�VNzR��p��&2��B$T�*��^m9�$y�PD1�4X���?��-���?����u�r �s����9�����F��8�{���+���f�ژ�)q�4\]0yZm�S��H��o�r#^%.y��Di4���	�}p��V���V�Û�¿��ў��{�S���Q�т���_n���7,�
�@��~�>lzm�U�%�]ޯ��<���Jz#)쏕����r�>���3��t#�&�>S	)��5t�O^�.�Ƶ8�U���`�`�.����X��Q��F��%��k�
�3%K/Aڋϊ�/�X�R�`Ӗ�J%��� ഺ�H�)F��OAD�v�A���*db�9�rM�<��:y��ś5L�ir3�&��E�X-Kl�p�r,;���?'[�{�ނ�/=t��,�p;�W���a6�)�}���
��2CP�j~ø�JB�?������b�_��qˁ������%�����D`�x��!�t��b�m��jRk4K�,��x��(]*Ӯ\5����q@�l���է0�|�u*v}k/�d��(ޱW��ዛ��L��,�V5^�I��ֈ2_	Gu����:y��
fu��{�	4d��A���D"�@G�W}K�u���Uo�M�s��Ik��M�̷�<]#H4��'�'�P�����0�d����-H%Z���V��\*�Sy�����;ޱ"�O��:\�>\����7�<���>�fy芔�����v�m�^�u�N�@���+�����a��[>�����VS��Ǉ��2�U8��3���i���� m*!n�07�ʱ��tG�z}tT�=
�{���B{&2r�a?_���8��*Yø?�E��8�k�o~
|�KV���j���,�WV@�|���|w�_Hq�*�]7�%>g��:����T[��!�����pڻ���A9��0�#�]�'��b�9J�y]�2mh�e6w��hǿ�v-�JXA�����8� g�O��L{*;�n���<���둉�O"�n�o��X��?Y�pw5���������Ԭq�v��|�-�e�D;~[���P�`-)��=�oAϋ_N��~�Ш0��?Di0?*�ߪqnpz�+'��%��p��b�7�5Y#6p�$<���vC�X��,(��?��-:�m�Q0�Ś����2T���\y1�h�O��Q�kL��J5w�'e&+&�7.��LY����O��3�7�n�3r@���o�N��q2����S���Ԩ!��w�L>��D�^�"U'�����F�,4�������,�|7���SY�b~��U�@Y��O�ޣ�](��U!�-kM�'�$+�����9�W�$����{��V��0�mR�{݃|r{D� 3�wZ�\��5L~�3��V!��(:�'�Q�[z��^K�l�MZK
qLC�˷ZU��B. K *�p�zӗ�B�%^�b��I@����d4�m��4��uTt�����Ș���ᑄ�x����Ѥ�hVe��Hs�\뢟��K�t����?����;��yF��޽�%�B��d��J�`{�QUa.;�A�h
��!���kف=���#�������@��e�a�6��C�>�B�鄰�'g��-���𵦟�J�#�S��d�v-|뀊�'Æ%&&�lgȯ%�o�5����-YK����%�-��0׍9Ԩ�S�~g�uXʉ����\Q�Y���c��@(�䄸��|�MS��W���3�F�][,����(4���zзɀ���7/S���[4(P�W_�h�&
]���̖ �y(x�G>������y�*W�U�:�*.�qp��RSd_P��0Hʪ�9�; %�4���	.BU��������)% ���b,�����+늟���(�A�cE�$�@�
�!���5U]���y���`�6zF�6!�Ć�* ��^�[�$�����H�Ih�-�8��7�n�!&]�|��++~5M6�OZ���J��Ė�������+�E���8�HS2����SM���{��i����bK���W�j]���&��`��5w�t�X֓�6�Q�.����9�!�f�i�B���s⽧���O���Eus���i��)]���p��W�g���'��=��6�C��1��FIq]��)G�G���@��`}H���>���)l��wr�KjX�+�_řL/L��B����o�2��O+��F�3??�6 ,�ZC�B1yo�wѺF+�Z@�Qt�r��t�x�D��-<PI?	�i���@��,[���/�Q��8�>uu=R����K.�R����Qjlo��t���S]@�Q�Ɋ��Ỻ(�/�2�E$X�x���׷�E�P)^s�O8Q��Q� D�=���i!�4z~�Վ˧uy�MQUO�q�&���lRQC��v�3� �G�(�zz����_Z����j��10������شXa��J�E���y0��Q�Y�)�d'�H�k|a��#���D_r~)
��(�{Jr%������M9��Б�BFa�w(1��ڮ�|��ش8� ��� �.t�ePǃ��c˅dܰZV
�k\լ�5C��V�g���c����fp����)I'Q~��KD钶͍�]�%=s�ط�
w	��945;S�@�P���-O`&�v�o�L@@�V�n�>Ӏ�F���?)Ϡ�	�J��XV��z"&৏�{��+�@�<|e�T�����l_�r����6"T���]A_�O��?���-��vή�91��G��)ó����f<ӟTV:4�t`:�����_�e���<��F�܆�@��F���6�ӂ#�����g���à�6������*��68vh�+U݆x��9{��2��vDv/?�O�o���6�G�W}Ų��[�����.���|����'`���n�� +�<	�r�CA=����{vq�gJ?��=п3�JI�ށ>�%�>���a� R΅�*­���v�Z�袲�v(����!4�yĬM�n���\�#���b	b&k�r�6�$�R����ڕ�aIg΄0m;DR�o�o�ͩAc�þ$7nF��S��<񖪫7��N�g�~/m�ig%x6i�e߿�g��V	���Q�dd������T/$�y��T���n�����}��#������$��`OۛO'�E�A�4���/�)��]A�^ �Y	�I	˨-���^��DVu���k2[�}%��U�Y����&�i�Z22Uvmb����E� �c�øQ\�뻯�.+XM��Y~�����Q%��RgD�/�O���Ԡj����?,�ͥ�bl����>S�^]���k5I�4sJi9��ri�HR{���,��u�zt�:B:�.���e����@d2G���
v���K�Wwy9�]����bk1�.Pqf_g;�m[�� %Wg��$�3�l�|�"���6ԡ�����]����
�"wM=E���fMN\�0�Gwm�R|��?�ƛ�row��Kޖ�]7�4���i��/���+��{h̳ߘ��6��p�a*�Sm��S��"�u"}a8���?��@Tj���w�M2�{��M+���)0�y�	� �&��!]_���c�)MU���c��R�<*,k�,�٬��*�m1ZV�$�w�q@M)O�`14Z��j��ԙ�|�q����`�� ���5����N��Y]=�RO���;,��A��%�F��v���W�sҰ�O$�^��7�ݡ�rYF$�F�0����1�".F3 ��K��M[_�ת��/� g��χ���fMJ��q/�/P���]��镢w5��K�^�*X��m;!I`nw?��[XKbT�=.�s�є��f��|lp�$�s��z�(��B�"�ep�}F{5 v۔uD	��w��š���cI��ߒ-��e�3�M NLb�qL��W�R~IJ��
�� �U�FӅ���ZTgR�=Lk��jå?{q�!�]s�_	X| w�JF�I�hƎ��v.>�����(^��En���j�*u0;#�v�W��O�_^���^3N��N3c �[L0�,���b�f��&k�Y�Ν���Yi����o%J��6��:�Or�ۖL&���L!y��w8����za�Yf<ڲ��"�2���/P��{m�8��}seV>�����D��B�C�6��ʁF��uZ5L����n�X��W<n�[m$i��V-c��� ���΁ԑ��Vp���l�O���oOA@G8���R�l��ۉm5��;�BB�SD���m�y�O�h��x�Ԭ�%wnP ����sk5Y��}��_����H)zV�\?Ô�s��盥�}��-=E�Ag��y��b�8H'�C���)�Q��U��"�0�S���&7h1��HU�z��7��=<*��,�xoUe�苯PC�Z�W���y�'��۽4\���5P����W�_Jx0x�/õ����ϱ�bt�L���Ǔ:��F'7�e��~}�cV��X(�c3هUG2AAV	65ϻ�&Ye��B�	
?��mq-�D��H�2�����*������`�t���@��)r���=C���N6O�·j�=q����0C�(��؝�lnaQ�<�lg�,{��)�+�����\���%kH�2�O{���$�o^G o�8J<0�v�N�2�y&S+O�MJ0�Z��l�>.@Ǘ�va��%k��-e���[x��>��΄������VZ��HnR ��K��%�rm�x��%$v.�����L�1�W$1�ե��K��^�+{� *a١5��!����Y�=��k;�m��*��1�{��E�*X�h,��ZOʕwxi1 ��� .*e� ֘zWԨ��+��������;u�)���KWk<35��+A��KvTv�n�K����o걽�ev���e�@�O�#��/�Au�/1V,mM��TF���Du�aC_��Q��ˑ���w�Չ@�;|��c�ݍ[
��4z�ߓ��)/`�@��i2]th���jwb��	�������DҀ�w����n�����{�n�ӆBꨛ�oo�ݼ��l�
�1܂��� (p0�ԯqquS�WC����	�R�E��A�����|p-|[�(�K���{��"�V�]F�!G|��¶Ŧ�����v��K��MpE�sE��o��Fi*�ɖ.#\�x#i�cx�;�t�T?j�����TO�|��z8u��+��l�75�1���!?��i�R�e{	
F��UL&D�	O�����w`�����'�MK^XO�=$ TE��c�(�����E�71�_�v~Q�/zv!Io�oƔ� ��>���Lig�����m��0Z�.�'�W�9Kd�b��#p�i\C$|����fv�0t(�K��V����������A�1VO8/kQ�u5���J-�p�J���ћ�ս�������!=�ay����@�)Q�Qh"��/�:^�����?舌2�6t�8]c��;^�8HZ@�Ps׎Ӵ���
w�r�j��sM�ί��w/�c�ڗx����� s��N.A�☻,���5�,`��W�ıg�$?`���)q��o��|�zõھ�!��ӝ��:g8�����/�����f��	�T%�ా��(��K^��U2����7���v�bgXL�lF܂X�^g��Rf��X�p�(=(p�4_�;N�i~�>|
����{I�f�Sr&����?G��OLFg(�47STR��3^�������O�ز��'�ʘ��,J&�s^��R�i��V/��O�~�[���3��|��k��˷�/<==2�6V.J��3�i5ȓ���� J�U�@s1�Ze_D?��k��������C�:y~3�������0=�����iy��t{X�UEe��3xnR�3R����l��͊���ل�-��6��;���N�ucz�Ry�j4�q�.e�%'Uev�ɓ�F��L����,A?�*~Ѽ�.JhY[���e���t�{
�jcϡL_,�o�r1E�TI���������(�e�������C��p��,h$Ȧ�
�2+�xC����@�&<���<�H�^�Տ�:@�x�3�Aw��0�E&�{���L
Ӳ~`��6(][��%0B'�T����[�Ĥ5�v��..)wN>Ð�;^��Cb[>�����Nr�6=X��+��d�1���N������ \̴ߓ5`�L6����\j�RB��άG��xw�1%��|��)�_)<jP`T�!�w}��R�ϕ,�]#Cqe�&�����=_1`ȉc�X�n�6ca�'�9Ě�
�����A���;�������&��Ԫ���(��W�rU:��k��0��޵Gz;/��f6)���B�[��M!��o���\�'6�`l�<[�����^��IA�D�a�s^�����aw�>�Yo#�'��M�S�����Q�FC{��o�ت��%�`��2y/����v>S�sNݦ®�~w�m��w>5'2�+�K��k��{������OfɜX�F�%S]���&_(�0J%�Hͧ�&M�j��d;Z��r��g���K���:�2}	�k6\V	%��sD8���^E)I�-����:�`L�M�\{ӻG��v�W�/ \���.�vY W�ԵM��QWG������nU56
ӭE9��n{�Nb�k��U�*��gO�;= ����e�C���S�>b�zEe��s��YԍdK�&�d�H���h�wm�ߝb'ό���V1�u<�\�� w�+�W��Mbv��l�D��=�mt^������o	�ƿ��aGy""����8���՝��/�y��8b`�tyU/
2�cqe�+ �9[@�G����^$?��2\��6�.��*�<�p��.�}r���� �H�������
�	(�A?7��ZLs=l2Z�ێ�m��$���Ƨ�R�a�4���}ݠ�~��%]��W�"�~yIZ!��b`�C��w���V��a�cG�3&h	e1�Q�;d:� 1�Q�I�0��I�����n]C�3��M�N��T����7�����>��7����ە֔4d����7���O<j6�ң��7�SQ�wzμ�hF[��O�m�ڞ �r���^��U�Ό���3X����<�ρK�q�a{$�'n��2询�N�F��֜`Q�c ����Ix��jk�;bژK����&�tH�.��7��?��o�k�:���w�P� �v�P]�jlh�G�yӪY��q��I�apמ=s����h���|�c�
�x��U����H�7����������,M-W��;r@�Y�X����E&�y�؎t����ʏq7,�ϡ ��������z����zϡt�ԇ�/s�(��}�1�J��1?��T�u��#�vB�����4��z)åZ��A2¦�UI!�5�V��`��aJ�"��<��<k<2We�W+c"�l�O�o
	��x�����O�](��8�g�7�\�x��A�Qf�l�݁�
��Ą�
���2E���W��'�e2Z�������*��?I(��5A:9	&S�Ț�&؂4�0� ��wa>P�/b��T{w{���OY�kXj��Ͷ���(�}���)@G���FK��}B!�����)��@i=�1#s�{� 6���n�"�6�6u�"����{��Pi���j?�kI��dze���A�|�^�8?�]Z���J�
R ��O���*��R(�A�g&v�5'�yP�-h9�oa��:�oн�=��X�8o����4~S���+�0Po�eL��l��p�o��$�����$w�)8p��M�M<58$B�|!�IM����b�y(ϛ��!�"�]m�&F�?�Hlz0twzD8I�iG[S�} �_h�o�C3w�C6��p��~�ο�����(}Op�� --?5�PE9���ob���8�����߯����Ч��� ��O�P��fG1�`�u���:0�)d�n�*Nfp��P\@]��
!:e����]hk׬�s�$��u�F�/�~�O�]c%��= е|���F���x�/�E.l;�����b��zK��EM�?>2�%d䁅�4���?CU�t���-��*B�S7,!����Yv"~:eڼ��{�M��Z5E�|RYx^U%�n�E�.��IN���|H��0�R�h���*���£�oy�k�p����`�-�wi)�f�F��x�����M�w��?ӿ�
�J<`��2llp�RM �x��b�����E�����y%>�R���C�2
4*9n~��P��`��������Tܽ�p�r]�F?9-�}
b+G����^�Մ
Y��A_�X<=*�.��H:�m�5�KBI�?���>�f�.�ɷ ޠ|f��i&�@sf�O�����[*y��F$\��ۗxre}J�Y���4/�EY1s����1"�u�J���F��&���#A��1O�\co��}���k��H?��|��M�Y���;�������i(��X}���ئ:��-�[\�"k�쇖&х������"���=�G4x�~��)�B`P��z&z:7}�zdB����$��90	�7�٥�4-��b�_�v���)i8���i��Y3Z0�bEQ��:вK��%��],'S�BV�ghd�����������.ȍI�I�D,�IA�>I�S;�s6��K�md�� ��_���'�Y�3��G=$�Ӳ�s�ĭv.r]�;�>e�!/��ǁE���j=F�1:!�h*��,��U0�]�
�I"�q���$��<u�"gԽ��oܘ�p��^额��Kc�!0�P~O2C��@�Ś�	���1��r4�/���(h@�3���E�7�w�M�����[��.��,��z��Jߴ��~͈~�4��ѹ��|�i���G��y�_��7_�.\C3���<ҍ�-ݸ�LZ���"~7�B�W�0��ӡ�*�c2㓸�b#u�������w@TdH��V3��׉� ��;�P�^�����bV�A���`GD#��Ij87��b;��׭��q�i��v����FHװb	�0���&��˥,~ve�( ���uӽ�$d�յ2��[�7�y��������b�x��@����k�a�l�#\��^kVZq2��
�;��y�"�k�6KȄ�-������1���T��tc~�8�m���i���
�*�ع,��,,�3]o�ү��p:��q3o�Ռ�Mۚogw��}{����^�?�c�ؼ���X��v媳��f2G�i�1��p ���Ҏ���w벎��M��P�|_�	@�r/��pE<��]\j6VRx�"m��nO������c�I��ǽ�Vb��ƪNl���D��%��ڛ��#~O1��(0���H��B�wħ� �����F�E�n1a��y	#���r�z��ק��ݶ�I�1Sع�� 7�y�PZ�&�Xr���j�97���YT��>z��߶ozgQ����Y���S�"7���v�	��MO�h�_�����1lk�s7��ߛ��4�0�W����;�!>z�D���Xl�PH��^�#��zp�؎�D�^fKJ:�TOH�C�H�w�����3p�@\�N	��}�WJc�^�R`�7&�A}�8����
�}�2��ɰ��&i���}��������*����{"Za��������Q;8�GTX��V��������4߀������p��tϐ����t'�p�d�v����[&���Ng���4Tԛ_%�|�����-�����ԉM�CQ��jPk\9�2J~w��U����Q�g�pP��{��;&V��熞�'9���y��`U�>�-�n��3.�(˻�z��[�}!<���&ß|9��� ���k"���a�4PӾن�p.��T��r6AwY�?�����8�2������P$�1����(Mfh����)7S� HH� ������k`�����@$�ь�r�Q�س)�T�:�k�t���[ͺ[��X�*��h6�_�ӤS�)٬U��bz�1x�u�,rR�F>��L"{�=N�������Ť���1�L�=WM@,�s�J�J�b�R\�?�3u����H�T�1֋u�\2A2a�𵩙�Q�p�'i��_Μ�I |�-i���&@������K�lLx@g��[̶>_R������^�.T�X]�	qn$-~���E2�I��#ųĥ��r�	,!@uV�S�$��u��馔�����n��okD3n��'�`�ĝ"�������zS�6,P��綡�9S(b�Uo[P[Z�=e�ijj������X�k��ϡ�	�P�|,��/��HE!�cp,�ts��h���5(J&#��Drl�~���9l �n��M�n���&c:���%=��<* vb{v���x	g�)��|���
2�m����f�ڕ�,TU���x��v7�5s��Y*^�&GL������o�ϰh�Y�H��G�zN��2�Ҿ�,�{��}�K�^�?���	�K���2�\�7�y%�a|��]r؋2G��ځ�g1�Q'C�b�w2��-��d�Di ��H6N�>�ǧr��9'�AF���ChZ>>��Uw����"ׯ�ŵ�,}=i<�c�)y�t��m�z'v��.�/����=j�V�ϳ�8Ӈ3d6Q��a�UQ�G��'�K�53I��[<fݎn��B�-31d������U�ĀZ`���8`���u�j:tɇ�Nl/����q@[��/�7�ϝ`�������уG��c�X��mh���8�d^�\�,$�)��b��`�>��yqL8�K' �Z�ƬT�&g�&���Tq!0���J��$FnT��i�tP�sȨ���F��4�)�;@I�� `k��k�]�[�E�1��_�p�	�/��N{��j��h��[;��%�P������ޠ��Ysj��WtD�����=NE[ ��̭�b��='B�R�	1�j_W[3��[)��I�^w
>�eF�qv�8�Y_���I(�EJ����C-ubi7�H��K1.^��rI%OJ�F�_�׳rX��^�-��N�8��At��<&E-<6���� /v8A���ӽ [�����_l6|�U|0��rXOP0�h�����\�rS��n<׳�4SPͣ��O8���5e������G�M<^ױ�����ѫ��c����Z!�Sk`�"dm�n�%�ŢO���	�0@�y�E�WM-��̇��J����Q���.G�|p I�p��u�b�Mڜ��
Z�K���Ŧ�����F����08�]0 �x\�\3�2p�E�� y������W]L�ʉ�-�p�
�]IMQ6�
�4��O�U��p���'A�T���$#7��-�lC�v� �	a�H�T��F��Qk&�=��@X)b���a~�����h��\f׋kf���o��-դ	�7"��N��(@k):%G�l5 ���W�z���\�
X&��fl�e��sE�W�jӿ�P�Pq��R�I/iB�\:���n�,; :w�@���RL�Q��ك6w%��P���WZ?iXoa��H9q����s[c��@�Q�_%�&yg�h3�	��+��>���m��ʯ �@K_&��r�;��j�i��C�d�����\�I��)�8_���P	U�!q�8*���{�:���{���σPMzs(�7+-0:R��%&��6����D���9�o�S� �����T�Xi�yڳ�7H~����_��1����י���뎜H��N	~��ԭ<��� )Ǹ�H�20D�*v��h(�����*N�l�>�"�ؑ�"�����3���Yz���U\u��1`�(a��ʥ��?e'[��&S��I��G��su��+P
�zrb4!b��'3���z�-Ƅc���nN���*�)�j%恸t����J!i5ɛ
Q��&ː���N�G/h�Nm����A��h�sSX�Q!ã��S���V����.�j��3�JĩMК4�����;�W�XV�Z#J='�qB�8ꈤ���i_M��XVA&�i�[��21;o͗�͘wy˪(?]"�iu��"�{j���τS�D���՛0{���QZ��Sz�X��P%�൭�}O��Q
]M��7���>��q	fi%��t�6�Na��N(Qi�������u�����>..��jӊ���G��~��iy��Yɳ����3ټ�b��o�CN,��s��Kv��L{p2��J�s��6�Q]�H�l=�L���t|������ �D�5@BK��w�J\4� Cn_�w�,��J���d�p2�+�9S��$
����T���$'�=�И�W�{{�.cy�Ż�
?��O6{�{����d�-,�A��#�g���=�#��1�� P�����!���è!��KT_�pihK*��b�D0 ��s-,>�̴p�r٬���:`�wXI����X��c>|~>�����Lx���a���֧!��p?�u�b����5�Ǌ��K�]���� j��J&;z�:J\�N��$D&̇��H�<�~W&VQ���vTq�	����=<�
D��[���p��̶'�Ƭ̅V-澙�.1��9	��O15@^M3�����T;��ۧW�v�@MF�'������+b�z��EZ:��!�#���&\�s:wՒ��p�_�-H,�\b�XQ6���V�}��"w�E��ɛ(�E�jf�!$��#W:=e�oz��r��r$��3&F$��I�pA��#[�WCt0�9��:�:�7�����i�T!��xݨ�8%Ř7^|�6j8���:��`k�P�2�Y�%v�1D�S��\�``���(KK5=K$t���n��2@�v���7�I����^�Y���R�'r�T�A��3Ax~��rp�dȺ�ǂ��'j�𺠉��E�#��M�Q7+����[�M,�nvX�%�c�^���c�8���x�H���m�1[�\5�X��]{����7������V{7=�"�@h����<����_�k�e�|��9f?�G��9�У����l�!R����di9?\�c,�S�:�j��{fKa-rz����[��luKB�97�4C"KY��ͽr�u��a��.:����$_�K�)?�}EW%=2�(դ_63X��w}���.� j����U��<_�ߚ�`�Q��f�7�Bn�^���B��o�!�`
qҡ�NڑF"I	��6��Gک�ꁰ��F����R�5��',}3;#{4�nK���x�{�;Pr�����⠒ܩ�0��G>�(��BPX0���ڧ"�ŷ,5��h$3h�<�	�)��r4�)~H89�R<�����¢��L�g@�4s�%��O&��S�@]�������3>��h0�OF��V�B������r���\Xe���x�yw��ruH�7����-�W�	4mXW��^�NC�jkL� ���<����I[.Ge0�֖� p��O��"�Q�v>}'{i	?�]�m@�F|u�_v���t>�����&\�k��H��xV[�N���~���a��2DZǔE��,oB��J<�	C��z#*�96N��~2�D�[e�#芢gl3�;�Ο���n����<�l�>�P;�v�Əo���p��"gQ�*�@�{�F�*O�	�=!j��Os�7.����)6uN�l�M�a��s�Z���*��O�HcL��݊7��0�韊'�9�8��N���w��ٍ���_� >o��.ZT�}1j&���4*B�~$��|0�ff��X���2e������caP�\E�V^��j}A���<r`�Y%rAbBr�"�\�[��a����+ 2Q�V3J#_�JLl�=�+F	��̈́(��U����s)	T��x�c+�a�]���oQ/��W/I3�b\���bY_�@2[��6Yϐ�e��YP"��� .��;k�[!��ƆX?q��T8_x�H�:1r^YKR�F��p~���I=��	���{�_��,�p�zt�K�J��˓J�~4²�Q(H
muP�u��(L����M�n3�B_'�W���Sې��	���EZ�,�^pU���Ku���D5��w '$��e��Omw�o�ig��]O{wA�<�2%M���iQ���vtR��&4���>��/��J=!�s���Y�դ��^��Ó��Q����Xx�����)|�k<�O������zM�Z9�c���k���;=�L?*��;�\�A"\M�t[�ӆNԎ�)I+��oV��waUYv�2���.>A��q�)8~q+BW��Ӻ�W��̤��\i�]wb�˖҇��R)���u�P��(�2�a���H���V�[ ��1WK�]孧?��Z.[�s�(�$�������lG`P9���t��}`G4.��
m��;B۬�I��:RΆQ�8��IM�$��ԡ�͡�2����ڐ�6I���-W&tʢM�M#�L�/�Vت��O-#����>��ʞ������{z�c�z���{jw|*'m���Ǚ�yk�&���T���,¼��iT=,^�P���

!�y�)���b��%�q� �]P�M^j~}8���	B�2�)�f$����{o�|U����4� �?�a�� 2����M#o�m+|�m{ړų?�\zɳL�m�V�2W��T.�`ru�˚� E�[�-aM�5.�����5OR};���(�&����B��WÄ�q�ǔK�����v���D�0�,��Oȭ�,�h�=��I��ۡy�ܭ)��¼����;2�I�����7ڍ5J�Iǜ�l�9�mD��7�-����7��	t]�j��a�[�[�J�ϊ�E��7M����~�j4���/��?�y[��EQ��F�3�^7U�ryu	�G��Ir.=9��[k�;�"nv�[����O�˲�![[]�YY���h��><
��S
���y��J��?��-�u��2L�쁡�r�CQ�Äʧ:�i�a��l}R��N���|�F&AM�ב���DS�p0�����@+� ՠ�N��3�E�5�}xe���=�J�����ڰ�c"�]��,)*h������W]���� �B)��W�����}f:v0��ѵ�0@*"���_9ʡ7@�Zʁ�t�=,����O��^9ŧ38q��X����C�G����K!׍a$� K��倄T|���P8�M��/FENR�V	��p���a�r�H)���עâ�*��LNiO��n�n�l��������X�%:���_Ƞ�������
�8O<��"v�����#��U�iw�s�-��HxC�[~e�~8�9�|��MHQ���6(U�� 8;Zh�B��¼�;�����?3tۺ���ws��8_�� ��~�4#���;�� s��w�r�b�;��zq�
L`1`�=�A�
}PS�ʤ!F�t@ݺDޥ��x�|
���f�n��e���7�bB�O����t�y�f�E��אM]u'�����.����#9�he�ɬ�T ����i�S��Oԡ��Wӱލ�����0\1���9)��2��4~l/M�^]�<�ԑ�AU��3e�Gƃ�x���C��fz�Ǘ�Ba�N����$���.3:[/����p>�{�`Ը��r �#j@��t��!�wA��j�Y�u�%P,;B�-���`�5s��Ǳ�k�4��X�r�Q�#�,�ȎP2r��0zRQ�p��Ir=h@N�#:��#{�����q�V3�XcN��:;�C��:A��Z���6j�A+����A�s�m�CN��e�,��N��F�'����l��]�����"S���q�7��	I���?�HHZ���O�9��Y8�����E#�^u���!irZ�]bl�ʠ�[Xl젲wGRnt1��cQR�����L�ׄ}}߸Υ���8k g�(�Z�HOC?o=!�&�X�o1�3/��"c�������
�y?37������dN����D��L�h�d��X����5x����U��A��.k�������R	����"Ɍ�(���pI�u*�i�oNo8�A&r�>�� ݂�7:Y+Y�@1<����?�jP�)v0p�N9ʏb�� ɏ��'%S���V��
Y`�D��\'@&��1�ݮ�<%8�b!Qt� ���(���d��3�/�+u1L^��Y�=��N)�2���57����w���U;QC����5��'f��Gk� ���c��Du����gV��y�'sg���ؒ�Y��A��3�vҌ��e��T�Jf�������_�SxY�n�-���ǿ�2X�3��L�x��u՗	�B�����3U%J=�ߝ�P�#Ee��i����%�A�V���%���`t�E�!�;�Bj\G~Q���?
B��yS��y�Û��Yk����|�*��ڼ�?8'�պ<G[,_N�Zu�0���}c�3�:hL��0����tA���Ǽ6ͼ$vl<s>J��J%��\��H�cB�&�R��:ۭj�%�,���^�#��P���}���?i! �qn������Z�Lo�Xl�<�5s�m㲯�	�j�,�^p��k;��`Q�������-����6�!�3������gOV����0�A�Q��,�Ki�]ya���Y��V���y��n+XGW���㡠b/�U�
<K�ӹ~avU���p޹e0�uiTM�%���D7���������W.®�s^�`�<��m��m�y����竧�O���7�����,�?�4v$]���C��A[g5�
́�	���c9JŐ�eHѩ�@?I����n!]������B���H֦�JI�u�_"�H3/Z�~��!+�E�>�Y:�$d
�l�Iz$�d�Hot����&(k/���x�fO���:�5�L�^"�x)A��$��ݙ�a���O�r4^�3%#']���I����Gi|̽w�!Lu%��o����Y�����H��aa(>��?|�x����G����;�w��+�A_mW�nG�J ���<�+�]oi_�JRp�=����� ��EZ���C�n��2 }�Ha�s�=r���}M���ʌ�J�c��
"[���7\g����GD��o3UԔRXH����-,?�Zw�Du��9���"g*�$/`�� �Q�!jn�}zn�-Hn\�����fV��J����^u��Gv`3}��Q����:��x�|�R���wW �Uv[�$&/�>�*�7Qo��e�p!O���G]������kZu��Z� S�?ظT�	}k&��k(���>Ic��xO��3�o7�v�5��_�3`�-�?�PI-�zq�+�ed���~�>�n	[ӌ�P��Md��q�t@�4���;,W,�0�s$5άNlc�pK�(6�g���"O�tf~9�h�H5�*�`gv��R����R��K4#���\d��iS��2��0�V{�9��ͿD=��Oi��� ��2]��_��r�;b}���8O�GXbZ���Һ�`��
��4Q��y
����&N���+b�PE�v��t\,s�E����!c��9�l�F @f�F� 5�������A7m1ۧo0�FRzV�)�h[�b��!��[�l�{]�!0RT��?�S>^]���qF�����D�j�@��Y���,�UDg����S2R_����ƴ�����j�k���㈷����=�Yh�B��9̵.3!Kd�n��:���Z\��Ӎ�d��gݺl�?�D��b�f��H>��\�_`�$�t��߽��������öա[USq�%�ӖO�ᡚfW��T�b�#8��͘����~Z>5_K�;����א2�����T���qT�y�=��!	Q�j���Y2HL����ܝ*�Tq��>@&��jaeD&�l��n�E0?ސ�d3,9�v	P6H>�]��>�XH��QA�Q�*�������
0ԇti~7�(�1W$�y�����;)ALP;�U}���?�BtmSމ��]�!��C0$?c�e�
BuҌ�����t����rQ�*lSp$d�)f���,���YO���pJtr�æA�¹PE2
���P	���s쑲�	OFL}v�^,�hh�H�Y���B�9MyL#�Q�bc?k�p��x6����
�@F��Y5������|��2��گ�ׇf��������^��v.�S��K�$T |�HZG;L��qv<��<�5׹r2{�0T�� |@���٤+�+���]$|��K�ߘ����e�S=�4D��jiL�;��3�^�-Ǆ:w0�KD�N4�H�c�}g����3g��45���J��+���pLD�+�Hּ��:��.Bj�kw�+��� 0M��źMp[}�:EVt�O�����%@���r.���f�|��N�fqɸ�LeV)T�.,.Yf�E	xœ�>|jz3�?���/���h��#е;��F_?&�&��KE��e���]τ���G�v�j��!"��m��!9���l�/��XH�
K����U���b_|j�G����Hvэ��Q�w�d1�SI��n�6��/'$��C�]E��u�L4Ȑ�W,�v���aI}��du��������Jc���1�#�z�5ќв=�	歞
��]Bj����)���!|�C�`�D�:8��~�I�.�J� o����R�T�U6E�Kq��Oq�EWa]Ѥ�t�?L?��gk�b��w�3:D$<(�~*T�C/+����ac����[�<��K3�D�r� 8�����"�Tt�H/�e�6	e���ɳ�J�4�z2�����"�ާ���YR `�f���O��N��J���6B�Т��x�F�����ԳI�'$W���ҁ�d\���VR�#��w���;��Rs����q���/pw����C���1%��?0ɒ�����B���M��Bu��]
��Q��D��6�� I�
Ԛ��F��l��6�s��\�8��6�S�t��[W�~��Rs��
����E,�"�P�� ���i���%�X�������*�=�!!Ie�w*\�$��#<���$<��ݛ�)��~4�8�)�w�i��<m�0ɓӢE=5&������ ���O��rg�bW�"p����AlЏx=��=�+$���\�����?�_69O��J/ur�t�v�A���K�b)��Ozw�$3����H�����Z�K{�7{ө��Y��|�
S,���dp,�])���1G��������tG��|=�QYJ�f�M9���9��s�8m��\Е<.��p!��(s亭��=��_�����?�]�lbA�HT ������N�'-;�F��rO�	q��1ı�Xؕ�W4Ţ��}eY�mù�=	���мu?�[t��Z�D�
�	0��ň��$��4ݷ���t7��|#�r��*5���gy�p8i��QxwY��+G�5?�������f!���Z����J��#�R��E'�P؄hTP��s׍:��6;�h��%S�����z���`�a�MY���U�?g�	�z*uȒ�/Y7��q�v>��o�mdŷ`���~R�{}_WU#{�(�]�ЖICv���jS��m56#��^�LW�����%��:��{V��t�xm��|�ŪP��b  F�&��&:�A�U�Ak2D_*ȟ�y�� Z�4���"}�#��eL���Ӥ��fH���\ė.�;���%�`�U��H�mn{9"'�6s��sE�f0�~Q�t�d���G�����A��S禴贊���.�<�2ᮙ�I*b/x)9��g��,ŋ��۽ɾ���6�P��p�V:��#]�j�ttA=�#,,�g�;�f�R������{��Z+��b�pg"2��*;j�~�f��%e�p�Q#o�1�q���f?�O��� K�CV��/�P�L�HVᄲBpX��/�Y�x�D�%4cc���Ψ�'��i�l�߼6�Y���ˁ�R���s�l�1�k��Y�P�� X��r��H��b�JB�]�EN����J��#�~6~{������s����=gTA}%���U���Z��L 5	C(�2�VM�6��>��F�xo��Ϭ��C��׽Ĥ�P�$�����/��)%(&s��Fj�^��4W0b�*�M������q�_��@��4�i��Ը.r��*[#Et��t"������ Ҫx��*�mw��)�5@�hla$����y��I�b�_(*�T��\�O2ڿw!N��z0��D�0S�UzV9{ȷYdOu��,2�)� ]�g��de�%�azZ�aLz��b�:;��ݵ�|I>,��:��h.㽎T-�� q14u����"U6�=Y�c�+G0Vn��P�[5˛�Px��> �s�B���b�Y���p�
採�����\Ӧ���������2��8o����B����i��z�e����8��+���kh)��z;d2�tl����S�������$G�9���c�����?x��C�9ٸ�C�We�p�؝��-�(�P,�����,-b����[��гc���ս��Ĺ�YY������ f,�t�M���+᤟p�qԵNڣ�X`\sԽ��-��Q1�d�L�/6b*���3��[��q���ޒ���~/:���vs�*������O�P�J�o�,��0W��E����@�I~�l>`T�ɽL���fq��`�D9T.�Z"�%���M8�2�i��G��Z���Pݿ\�w_[�����ӿ)���UY��W⿟,�M�Q��] cv�$�!{y�e"���/�}~�Q�8�(����o2��^WG����Q�b���N�vvWn��GԂ5A"���^�FA�_bV<~茫�_��=H�b��X���U|Ya;H���sNZ����G�vj�($0��P�]@O�/W�Vf��M�Xu����йyR29f�L��+NW/���8�eY�؊�̚pv ���(�tُTQ�nd-
���gRL�j���>����:�Х��D��hM�C0��M�b ����c����nT��ڸ�'�q2:��N������v#�ރ������ݻxz?w"m�VY2��I��e֥@O��M���=<a���-��e��٪�yru�ޗ�>�`�@G�q<����˰]����D&�7�W1��w�ѓI!�_��]E��d�o w�w���m �(� 
:�T��N;�v����xK|�����dTy��Wu�s�!�y���B+�)�>B~���!�U�$���33���k�P>Nho�[6�~f}*��ocC�]��VC�K_�~/�i�1��CjAUq�7�*.n{R�O�ږ*.��ᮡf�ȍ�;Oy>��P\����?���S*`��g;�r�$;яZv��O͹���� u�E��yӨ���d���[+��P��0�H�0��lB��J榐.׆S>�}mB�Y�Κ���?@<�����[���yo�]�]��<YR�$<6�_�asd�"EL��
�^�!|��Y�yZ~��y�"�9�˾�U��{�}�}ڢ���&�v����K���� K����YOAi�?g��q�@�y%b��hP_�$|ό �K��dt��/\�;H$I�пL~}:g!]ŵt�z�r�K��,�5Ϳ�ΪS�JD�:Ufig�O�}\9�NgQ��6�~B�_Ŷr���G,���$�*P?��q��A�;,.���չ)h�o"�M�^c �I؟�`�FϜZ��m.�@ge� Cׇ�4e���-7��l ��<���T�c����#-�U��>|�����v�W� �n!8���'	�{�G�Uť��e�-�깘��R��e�F�L3P��<}W��H��Z�I�z����Z٫�(�[a�o�H~b��-�3���f����^(��8�ԓ,��H�_�� o�=T�\���%�ĥ�V$ �@��e���ѳ2z��,�5s�L�[$Χ��"S�Q�� �wIB�� ϔ��-�݃`��>��M}�|�0��f˳oTF,����è�0|��z����0ٺ��*����ww�[[�&�׈�6��4��յF���=�d�s��4|{[�h�莣��/�Ji�R��yi��D����T`�X˕G+�iC�VD���]u�{8�4|.�*�f�q2x�'NL��T�q��G�$:�)D��|cn��o;+�C� �PO�uH�a�Y;��1�~�3���}�
%���t����_�0�cXH��\�\vA�x�ɮm��Dg��"�VQRTx�	U��*F���Vh�o���%t|�n�y��i������%��zɌ�>b���IǗ��ͮ{W�cE�[|�)��s�5����?�k38_�ǥc�ٝ���|�2�K檒،1ms(ǎI���(�&1SMP&��������y���\mar�Su��M��yx��LHK���
�^��k�zm�caϐ�nƸ}��W����[w�����t��:�.j�F٭��&`�����&�w��v1iD��x)()�ۀkI���ge����2��U#X��C<�ԯ ����_��*'��9,��������;3ס�r7���邗	���G��:ZMv��'!���$��w���e�+�u��m���u��i��GIB�w�c��A���z�Yj����=WP<ȍdǒ���pҀ�)_,
���k��K?��l�4���L��f.8E�N�G�>
e3��!��#Q	�k�&m�S}����'b��pc����1,sRwX�{�Գ���{;�u�<��+��#Ao�S�����Lr6�����Y�>��,2��:�]j5��&����v{4���� >۫�j+<�M�e�]�b�.QW����W[�Y�i���SF����R=� %cM��������yE4N\pi���]n?<H�r=�I����to�o���\�,Ǯ��z�NuC�2���S��E�Y��I�Q$�t˕�ұ�oG�Uob� �2�O�k����l. 
�WY� 5����a�B������]
\�g�9,S�K��\h�Nw2gVas�8,q�/XPKm��F����j[�_҈]�>W�j>P�$��$���?	p��9�ߓ�^L��F*�_��X�(6�iJ��A���)���"�m>�O$C�/tJ;G@�{I�x6"��B�8�jC���<�e����4�h^���Jx���a�uiЗ����s/����Ӷ��mgl#����N0�`��
ġ�/�i ;=>B������0��Kk�oI%+�!x��Sr��-_�D"��;o��OYh�Q)�ӣ���_��� ��ٴ��1��)��A9Xmݳ��2�^ѽ�����N�B=�[[p�lƻ��[,,!�v�K�i�d��!�?�,8<ġI7��ea��ur�{��fM0�X ����m�*J(K�J,�S���]>�z�~��C����K΄#f,�2�vp=�>o���B��N`����K����7�i���Am�	B�E�D�����@CM���ݪ��]��M�c��^�7���`��}P}̩�-��8\� H�����e"e�+����g
����M���n�^l|�����~��T}�8���a�N��q˄�L',��ՒA*κ���J�#���E	ԻQO f�jԄ��2�^��c���\;��= %�a�t	�Q5�����T��[�#�S+v�*2�	�8�1������R���S�;��"m�u�����H&8 #]�Ѝ�����2,�Ľ����=���^�;�)���D�,s����R��Ϣ�b������pmj�l��nͤ�k6�=����S�0��&m�<R���z����6�\YT L�b�v�b�B(ן>�J;��Sl��z�����at�c��	���Ɏ<���ni��OU��#lw�9r�吥8r�3eۅ,b��msM\�4ŕ]�sA���·Sr)IyHރ�T�[���`�h�

i	��
��.�����VzЍ�Q�0�~0k��{qwRNJ�	��|H�8G��yO��Z����yU����j�K�|�J����0��s8YM��o3���XގM�!�Q�
,B6�A>��˻�����9�?f�{��s��4������e΍=��zu�RXg�{���
���i��"3�8���T�iSµH��`�6�йK$a3K�
Na���R�7�!�pT�p�P(���Wrb\&U�S)AV��
7 ��)Ud�ʖ�ۓ�t�I�]�(%[XC�r�/l.͡W�����_�c8�����-@��X���,�pI=��0�����ӝ���V�YFo� ��K:�3Y��`*�U�� 9��nGd����0SX@��&�rzZ6K��χ	H��I�������w!�z�q�_���!W[���z-Y�:'��O�z��D�����:�#:X�R��Ai�
���8Z�����UE �#Y�jT���~�{�1�����:�Y�o-0]Mr=L�����q���ͧ�<ݦ8�t{���&i���c)WN�a'��j�!�z3��AЬ��jT�����]��0���=�n��6�f2(�#E����0�~���Kc����bC=y�j�R�N�;qaؽ��(�()w3ң���r)35�.18KB��ʿ|V�g�"���-���ǖԩ�ݧ0=�5Ȧ��c��Y�l���Ϲ)���T.���ֻ��o�R�n��� ;y� ̯}�p*� 驍���^�h��=磡*���|~�"q@>S'%������F�᜜����֤�H�i�g�l��i�+�1Ȉ3#��C�
��Aר%�rydc�f����iR��|AZ1�-��������H�O�O>3;�]�'_
>$�`�f�r��(z�v+�x��&+�7N�8�?$��:�3k��<�td�\�&�^��	3�*B�}���¤	�~�'*��/�X6�_�08����N��*ڍ����K`l'B(�����y@���~��}�$L��!�K�9�j9�;�]�0�=x�^�e^�`�+P"I��\r����J�C�6���R���m͸< /�{mm�5��^�^�u.��@�u�H�Z����;JV	�h��&N�k�V0$���܇���#�q3�_%-��Z/| 	��( ���Z��ԞI��<D�'�:�����BX��N'���&,槭'��R��\H�|Ε�D�w�m�ns�:ކ
d��Ecz\K	]a�f���da+P���������#ɉ�1��!�-a�]C�����"������M��Q��/?�A��(u�t��0�g���?o�u�<�Gof
�Zպ>��Y�J�D�?�ł(�_��~MRתZ�\(��������6g�r�b�,��}�$ғ�_0�}�4A��:	���6èL7޻���J$��y�o?c�y�K�kw*'��N0�:X�y��bvt#�<���n8�½�9��A������:��MԀ,�4~�LQ�{� 2���#�{��;C�(U#��'c�$�%W!�=�#m{�w�
{�s��D�j��` ׃�v-��J<
 +�%�בPf���yѾ��{���q��@�Pvݵ|�㽂�{̇�x���ޜ��U�CeDb:�Z��C�ȏ0�kc���7D��$���E3m�9|���\n�t�I�A< 3��T���Xo!��sJ�ٶl�%G��F4�J�3���r���}<��q����K��y������DTjr�:�3`�b!�ji5 6�`6���@�XxͅB5�zg!G�- �xy���e���Ď��[ 1�~�f0�՝iGCЄ��g.�)���4�
�ʃR��k�{�#�@�����O��w0��I5Z`���^��c��I,��==%Sq���6�`�(mmʫ��:��R�k�����1�+�4�Y������1>fd����&�7J$$���[���UX��Cv%N��Ѻ2�(d��Y�/M�	:��it�ԋ|jQ��\�gZ{>=���(�����s�n��	�j(���I{֙��|���h���M<�_?\�.��g9k=���-�/E�����1"O���w!��M��]���N���ҽX���X�Zf�uW8�f��i�a��ֽO�%�n=�?{k@�c����Ҫ�dŬ �_9;�R���|Y	��J��P!��u �\)��F7T����p�ۺ�0�a�Q3�N̂��i�Sy�3�A�$9 ��}5&���Kn���E�E	���c��EHKB��9&����mܮ�p+T��T\NU��H��ː�|�%A1R��P`���'�bLN��	~ [��l6"���+��[�"e��Q�ƚ�-
������--�~[�Ζc�g:�{}r�2:\�}Dǖŝj�.Ts��� ���&�(���Y����U�p�̢ǭG�'J�?�ú�G���4�N��h��mȴ�[�x/�Ѓ�JÎ�r��3�{�E���W٧��J��>ۨQe@�O?5�=��{#.a��iG�c^�]��D+����ѣ{b�X�u;>O�\��\e�_�Uǟ*-U3�{��kpS�ֶa�]�\y�_~*y��oE�U�	�*���5��2�΀,��!�`����,e*�֑)ܦ��6i�O4�N�#}��O�ʱz����κ�j�t�wq=�����?"|#˺q%�8wګ�W؇���M�	Hl�MxC�	]�N�>���a>�
������_���N>��9uw\�IJ��;oYlh���@	���C�,��h[�]���t��م��!$5�6$yȢgN��6�N[�2W�0O�L�?�~ga��ّ�����؆��?�j��������K����'E�~�,���|�����<�i�����)E�TX.�����M{n�y1	�a��nQ���Z�.���Y���leZ��8�[Y�|B,P">%�jj�|�~R$z<�9ln������h���������/�G�0�FxXk�e��nްQ��x �*�P~=��'��[�,N1I��Lt57���ϲ�x}��Q;�o�mԀM�)p���!�O��~��'(C�B�:]kPr2]��AhC]��;#�q٨�w�)-�?��⼕PP5=*j�P���ֹ���I)�R��\({3n!�����-{��.��Z|Y������N�t�Xe��Җ�߀��L���|��hA�7���Ƽ ۨ���\�ҙ&:�!�N�aeKq�M���|/�	����-}�(�}�}Lu�_��s�\[ !v�$���RK�������e�i����o����-����*
X��;~�86�m��$u8\���$xu�"�/*j���_`K���cބEE�Θ�&��6aF�%�.���5} ���i�l�3*W��^8d�gp���S��^�r1���c��]�&��Λ�E�ADU
%�����x��Ĥ�dH��d�0}��>�)�k�q?X�z>�/k�h~+� ��rr�4��pwc
6�Z��7N�2��ٴ��r-͢Y��2p[p&��Hh��T`p׎��ȹvח�!�^����Gi;.~a�'庒�Z,_�Uc���ے��޵u����b�8�<�v�/�T-��;6-=�O5��!/�������6��y���S�&�
�� �O�_�'ӇN>�~�����������0և�1�A����P���p���m���S�iO`�6�XG׌���c��VCN��w��Մ<i��n��;FJ�a�=U�9C	<9Լ�yұ�����`+��⤨��x��T���k�;�SQګ8O�Xu�2�2��)�6�4�� �?U���jJ���e�_�=^�V@���JEk �N����鏣R0��i~���p3��>����V��6t8[ѣ�t�OAS�u���C�S*4��Hz0�Z���@�܄ �%�x��N# ԳGz	�L;����SV�v�P#��4͘�G��8�X�$k��>؟+d��Q�) 6�����J�A����V�6y�gQ���U�~�@�mN��&&��\���� �ж��dm��6�A��Uy|S���{�8*���ȃyت�!x&���x�����K�lt��y�<ۆ&h8�
�V������/�������sv
g�h��%����Fh�u�J��-ǡGMuHؚ��;-5(㤍	�Wf�2�õŦ ՍbL���fS����Ѹv;2tH[[cz�z���
$��&�e����N� .p���4v7��ŭ&u�v���3�Z�j�p\�`2V��jj���X{��⣇GY@�g/�1���`�	R���΃Q.����.Q���ٰ��cV��� /y���2TM��B���<�x"_��AoO��X%-ӂrFw���[�����L��&� ���E��g�!�vj,��$Ђ�/����@�3q�b��[�g��lJ}�^�v��E@�喱��y�a�w��~�����9�W�R��������G���ɋ��Bmۏb 4;����hҜ��X��z0��溮X
ZI��N*�]�W�8G���ة�J��N�;O�d�HW' ����
��m�G��B�c��P5[BT�_J��TW�ے<	�ڎ0����	O�\c��la�"@���ov�k�m�d�U��.��+�{�[^Xݶ;-��?�^];�p��d1��	�Bq�<vUNk2���r��p[Ɉ���ز�8�HUf�+��'�\K�5e\j�C�d�Y|���B."^S+I'��}mN��2���Fop�r�N�H33D�7-����\wcNC��US��Y��^�&}z��C�݆QY���{���f��3�9�@U�7��n~+��I�,����JW�d8Ba��]�	-���*�,�N��d�%=d��u�:��eCV�^���W[!�:6v��J�����9L܃?3?I.	M%�4B��rw���ϡ���E��/����w�T�B��{V\�%���pzw�#XJ�0�m�o�!9#n�PB�%�I�j1K����
猋u~�^T��u& \��D�nG�^z�K���ON���#(�L�!&U0ɂl�cs�Pz8�*������N����p�e���ՔZd)-X�Eۤ��*٨ U��y~�,�z������/�	���
�Zy*�:U�<H/��;LY�Ɩ?s?�T�Gg�k(~���t~�Vʧ4���+� ɟ:��nv�����V"61V� ������'��.ؤ�#��~F,%S��h��ZJM�M5�YDnp��T�Qn��uC�����#���j��ؿE��֬0�e��t�A,�����3#�@C$9�o�B��r��5ؐ�>�I�G!���T|p���"��s�.�����;��x}\�C�(�lV�趌�<v���_>�M��ϡ�ˇG�v������J�7C�X]�d�Մ5�X�`e�����ܒھ��2�-m��U�~�V�*8�BLf���,g�,���]9��t���ue9��8��5N�(r�3���9r����u�����PJ��Mʊ���|��'k/�@&����#��}�:tHa���G9�r�M�-�b{���AߊB&
�T����sC��O��Q�����Q�Zv�����:O=|��{����Z��
p���������3/��/�UG6L�^/� ��.�x���q��	+�2�@�b6���Z���+��U�;�h��|Ôleȩ�~;�6��9\0Ml�Q��t�ݔ߃���@\� �mx.[��/|H��M��^���wA�T�-"!��@2E���g^Z�Z�-.v�΅5�vל��\VP{��:h"�x�a(�4p��󤞳�Q5�S��W���B��7��.-�$҃�$�m����Cz�>L�q�S���<�4��a���S
`*ihSꅅa3����O�ZY�rl���C,�}���n�
��m�����0}3��Ņ��`��r��y�g��p�zA�&_C��t�Q
��a?D�]ޞ�(��Í�� �ו8�0�pLG�H�3�_��_E8S9�[�0+i�&(�p��� �!50�M���j��'1�q�=[O"��5�?�����_��o�3�"�4�i�%c���TQOj�dm�K����~8Sj��kT#����[}��ƈS'5�j��|z��wXm�G~8RU|{,���&+�G�z��V,э�._m&v����k�z>��$�.4��s�G��d�=��>��g@���VyY��G�|"\w}>�6�"l��ؠ�,{��mR �H!���q"�24/�VXp{�B�U�ĳ#`5���Y�)zn=�Y���G	��{~�r���	�Y�'���Fl=2ߨ��3vF|��`���M�u���>\FC]i�)�}���~~���'� ��ι�|)$���{���`��e8���gܢz|,,@f9�l9��Rhz�R���~���qL��%n��F�?���o������k�bq�P]�^|(�-I�]����$a�q�l@̲��U�0݁����k����V����~���5V��n&���=L�K�������O���
�G��1�V)� ���������K!��܂�K@��pi-���)p��lh�)g05�j(A�Y�*
_�����H���}�}�~~������T�	��W��x
n���������	!��E���/��;����h�r�����$U����5��6@�h&��� �J��;9����ld���B��,�֩Swv������E�㣢et��d��a���7V�~Tɝ?o{G���yZ�;�����N�Y�����{E�=͎�<�G2��Vb�R�fY]�i�{��Qh�>[쎺��x��׋�R��f������w'a4d"D>E�(���w>��W96qۑ�S��i�f���pC�}���(�Q1=NN�/J���CiPO2X�ү5$w��?%�yD����uS�D]��3��mȗ~��9Y[	�ln���Ɠ�9c�P`;����խ� CR��Dc�FZ�^�?[���ѿ2]4H�R d�MD�M�*��C��VO����;��C�/Q.-�2s>G�Q�Y�q"w2��ɑ�Kn��I'��i�aOj�j��4���f��d9���֮̋R7k�2\N��8b-�
�,���ӆV�V�ȫ�gT�σq뼓�l�M'��-W�43�.���JA~�R�M���%<�k$��\��dKƯ�,���8h��ô&�Z/�ڤd��U
h��������wE���\��5�{���S���v�_�F�W
��䢐�	u���[��]�1����8j(�8ȧZGp���V�Xr߸\�>_��O�?���*^�z���P-��
��V:,����D�p�.NW�R%ɦ������OOvov?����9XG��W� �D^RJ�����$� �4�e��C���t_ݡ��-;?o���/>�E���D�+��Y����Et�M��&���d���yM���}�,e�Hq;` ����v��_�3�.���ԉ��==��9�����d�ِ��/i���m��&U\R��5��u��+�����'�uT�Ii�ʅ�Ciez��^b�r���u[�qL9J�'�5`�D��I� ��P��m��w|r�!�� �V�'3(� ���
��hVAiy�o��,(B�}�ݮ����kROw�q~&�MjG8���w[�@�ҋ�5~L_X@�<ֿ�G�\[�P������i��?��: 0��Z���X;|��f*��N����pfŢ*eꋳTk�zO��������X�i7g��(��!� X�R���F�~��}��NT/ʢ��!��x�&.sR6H���7�Q�4�٭'�@i��Rʡ{��uft���=�c �3�����Ĉ\ ���L�Rۇ���]���S%���{ݍ�����s����.x���Ե�*��5ړ;"W1���l�Q|�D�XG�6
���ܷ���:��\���rH�ֿ�17S�_C��UT�S�찂a����f���uqb� �Oa�F��%�����h�g/�l�0��#�;��.ͽ���z1�)��ܘ��r��(�,�U0�¼7�������gdq>:� �Fz��I,��$�
�瞘�j,��ި���\C��>=g(����)�:�r��
P�?C�̶�>��9�3�k�E�mol�S�k�J1�lJ�wGC>��ۏ��B�FN�&yܱ<i��9UD�H���ݮ*K ����F�A�|��N�1[�J������T����?f,�"��Bg��o;�'Z�����í�w���9���}�'@7�p�9��3��C�vj�0Qw�t���@�\��AƆw!�Y<\-�(\��Q�͊	-E7T�͢����?��m�e|�0�3���!VS^���S�-�$D�	ӣh�^O &�����e��UNcE��a��#Q)
�.��L�pln�ߙ��Iq��G�q��X.���˰�,]�p�yR�G'�B�3zD�ӎ�Ġ$w$H�9��ލ���	CH�o��,��)d!��C�l`/�:��@�ݝ2�A-!8�Yt�� Vx8���Ns�k��TIȚƳ�����`�ɲ8u0�p"J~�,̤�_�W]M �o�I�]_<J+6�\p��<�P��ɳ��l|��p�܁6pSf��;�S��k�E�*��|�XhD5���:}����(awA�Z�a8ˠі뷕����h������Y��y4�M.�]�B����>aI��7�
Hf��{	���ԩ�r�oQ�q�f��k{?5�3������|4ry��o��(��m�a-�Hh����>sq���T"/f��y���*`����0d�	iD�	�7��&X}��'y�쩷s�`K���4��*�%��{$�����\On�� ��tB�uH��b��i�Q�&����FA:��g��Ǿ��?�fNa>&�1�:DP/�mmE[�|�B�b�P�o�����]���mK��Ey'���'�kREl�s���F��������ag��:�PML�}�VIUD�c��8�[��8͗i". �]��o���<��0�~(�D��O_����[��s�1�Y�E��qM�4��@��P���qs����S���P�������O���b|�ذPي�:y4C�H%|i�[[��	��봰C�E �
��:8'��=�4���>�|��B1ķO	[x��Y��As��>DWNX���j��+���)�?3�*M])�q�3�ݟu�J��A��K����S��g�z nԼH�D� �TM���'���؈pU;�{�7�;Mښ����l%Ã�P��K�ʾQE6��3�L�������l��I#��T�i���jP3�2���������[>����KX_�=���7sMō�B�@�;3�ylhU�<k���5�Y�����R�J|�<��K��-�ָ��N2�o�t,��:�O�)���ٍ�wǍ�u�k��G*=�5ʃ�!�k(E����{�d���Eo��e��M��ߣM#�C�����h>�䦔x�-��5���T��ԧT/�[ǥ�yW�U6W���/���q�f΁?���n+u�Qm3c/^�J'�5�����ӳ��5�=�&����54vm׽侀ObλL�/6.��f}�8�L�	S��;t����?a+.*�+[�4�mLp�g��Ӳ�3�l��J�<F��d4���+�{h��lp�m����~���E܋�|�56Y�����q��-T�Tʒ*�t����t\YJ2�� 	�1@M�Y����ak�p���d�R�6w$RdI�͍kBN��d��	�RE�2H�Od��2l�Ԟ�k�*��� 
�47�&��E����
sB6{��g��$���e۬@�zi�SH-!�����3[uH�W?ݨE٢���r�t���Nӹͺ�������8��J9��s�@Y!k�kfǿհ���ewX5�x�0����\�1���Th��GT������_h.<�~ub-R���*�a�_�`3 ����V5���@+�]�|cL�6���h�F!�����5S#X��x+Γ�wG?�cc��7Eb��y 4`Qc������C)e�ePr�ul�0�r�v���!��9�c�4�+J_�B��ft�$�o�!��]Y��ٙ�E�i~���!pr�R+Wp��k����q����NA�����vTu�U�|v_�S^R&�W��=��Q�!�T��b����"z��lA���cJyre嵐���?��/���kh�ԐW��b�D���P��%lT}����n�x�� �ë�+B��
�b�f�*dP5��ſ�a���K���5�=����ɺi <�DӇ����q*x���u�Z^�U�̔^0� �����Xj1�<2��˫)D��C��T�w��<q4��?���)���E�k��j��|/ꁎ�� ������Ʒ��Erl�[�]�D_	��3H[&���%oӻ���b�[�A�n�߱��zٰ����P;��H�)�S��T��?N������]I��/��Z�?*'a�ڞ����b|����P�>J�Od����(�x�5 �-�U��B��-%��!!l�k�M��#W���Ʉ@]EK{M��q�fV��6��Z���D������,^6|f5���ݵ&�ol`�f�~{Ex����n�6e�e��]^���Zғ(��Z�{�g,wS �S#0JR[ыO2*x�^�wc�������ԑ�*�N��>H�����بX�	j�`�o���#�r��7�\�1�vs���M	g�E�����	��.@7���!����a;5.cZ����TI2R�́���~�d�R��uP���#r�h���u��Q:�k ����{�w�|*3�	yH=��~�_H6�/+5sH7����a`��'�4kr���C�\�q ݾ��y�@�����%"�̟��N�G]��am�j���*�<Jϗ�I����o��o��l�u�mLdXG l�A������Su�����7~	�j���/+��D:!� �
Ԫ��P]�#%��Қ- G�����
��S6s�� 	L�2��~�>�z3Nȷ[�xfeW�&����Lj�m�*�CK�@��8tI;��>4H���W\�8g�͛�Ep!XIW�H��$h�El�d�_sS#/p�K�4by�t/�i���(Iɗ���J�N��| *��F��Z�&(�mD�;E�c�͊[�IZ��A�U�,1�Z�76�����S�= 0����
���� �Z�'>ra����2��������ϰ{P��Qs��i{~JV�]Gd��ՖJ*��\�7R�M�c���k�&��i.�����R��q�	D��x�����JfV�)�d�<�^��r��$ۇ�{ڋ/<�N.= -�B	>�����hڭ�GL�<+}��zYEvw/�)gU�yi�Q*7�b��G��K�crP����{�n������1�J��"U�C�ƾ��j]}wwU��-�l�ݩ�uE]F,{�
�7w��x�yV�����f�}@�&Qcf�혪����)����[/3.Z���s���Nl�������Z`>u�m:��s����[��b�\���.e(�ZI�b�a @��3\��p�4{��U}݂W�]�7!<��ӂX0A�u�Zi�}:B��@�Jz�3�i�d�͘���J�WEzyKªh��wE�>�R����1[?�#���������ŭ���R �3�&�:�˻g�����3s�-�i]ތ�T��5�rjc�"u.�+cz98t)Z1��X�O�w�����YfǺI3d ���ѳl"�}���"AH�e)9B���	ש�	C���u ��=�J_�~��|�v�����5��~;Z�G�����W&�ډA}����H����1K� z`��c�F������4�����q<�/���e�՗ԩ��6t7��c"���<0��R'va��4�M-wİA�MaU)�gbRU���̇6ВtS*�O��ZM����fs�q+�@4�K݈Ĕ8�&�=����s�����g���z4�y>�]z�m��b�?�2-WI�DOAOe�n�>j�h�����n��=�"(K�|YZ�`���k�%�1-v��_ׅ�l'g��`z�� 	�klPkH"c&�.rW�m0)�g�S��&&�n��T/���Z������4��눬9�|p7g'�ӝ	� �4|���������l���7ְ!��x����5�Fq۾BM A��`+J��"l�wM���*���
uV��Ï�c�����szV
NHFʠx�S4�Pg��QV'q]\�Ȇ�	�-��{����2G��)Zk�/�؇�o�R\��l��㎌53�F�d����������c�Q)��+`or�<-ʳ��{���~g��*��/�0B`W|��j�¬��uo
7���DJ��G��_���
$��x�uXŘ^�B����"�)��0y9�PlyE�K��Iw�J�򓎦�-P �<!	}�ZU�����y�.�<��> �l?�w}�HD�ndi��5=�H3]�]/kC�M�-@���:�2�Aǃ���ah�(�}Ш$��I�a��p��AJ�H�f~�5���+fd#�� �����^�������D� %7'��#H�*R�ڵ���ք�r�">l����ү6n��m��,�f~$�[�;�d3�ʏ��ѳ���ٓX$e1ӻ�^��7�nF���=#�[UD��|VpL�ۆ�Je_7�bf�����M�4%�'L"<;��K�<a���9)<��PX�b�1l[2O#},7u�=������C��d������%�5�|��u����O� ��ҋ!�	6y�f��$����N���Da8&w�r���or�6�����@�WӀR���ɻ�l���P{7�AG���� �ռ+7~J
ַ���[ !����4tZ���|O�6zDU��`�vS�QtA�@%���n�;j�{~�8��d.]G$���!���� �|�t�a��f�x���9� �?��8ө�|�s�����(��J�Y���r�m�Oa��XV�\�ʉKM���b� �z��3
��z��(aw�U7r���l�f�=��=�xGrv��Ez.\EyNrlD��P�OB-�h�t�}au7�b�.JQ �=�P��ģ�ãf���W^��A�Xl�Z�q	���Ɏ��: �'��Ox'i#�=�c�3|)�a��r�x�ӛO����6+-mwA�_�rD"�N��)��h'o���m�Zt�sԶ����z�A��G�r;SS�ڽ4Ǿ�pnЕ�[J>����V���t����A�bЕ��)����?V�@fW�~����lgϞ���x��4�f(��U%�~j�'�Y�k�c�g��*��7|5������������l{��vd�Õ ����wy�N�;&�P��S�w�O��&^���Kܵ���]�#"d���xU���YIL_9%XJ� _�xt����^*p����#���E
���+[[�B�:��&�{�pwѮ��a|�ߜ���N��ys������R�ІGnJ���0��x�Sq���v_Ţj�� _����^����<O�i~��e�x����n��	T��.یn��Um)�(��ݳ�W�H_��qk�4��]͐�+�����հix0`6;�5^����s{�_�לm_.�{�5��3[��j���	� ,�����[�R�{&��g�xP���_x&�P�3U�y�����Jj@��%�`}D���.m+Q�v������BX���a�S���Y����ԡDF�9
���1C�Ao���k�>-Lej��E张�7=3D`�p�2������;���bM�
"N�9>
Dñ ��e�&]$��@���?X:��F��|�DGњzeB���jy����82#�� uK�Fr}��V���-A�z���|	��!�H��b���]�N��D���,wG�Ģd(�ӝ1'2�xE���>�AR�J�e�^��3KN�;�c"E�Ĕ:Kȣ���%[[���|{[H�o?*��]e�Pq�S1�9U���B�~�<�V"�͇&R��js�����	���\~z�xᕌΒ�t�饊*��3��� �@%����؜b�.�L;�PV�+�j�V���;���(�茲�1m�ެ��D�.rm���[�����}�|��o/��n&d�x2��'���˲�f�M!ރPT���U��x�N�5a����i�����Ш�\��Ư0��UhAS38@��N�7:k]|���*WM
� I�)���Mu���9X��3�ֈ'\��CU_������F۬x����Ä�����9 *�k|�>��-0\W�D�D�r�v�e����l@��* �������a&Xd����}h�x����t�(��^��1P��Y&Ɨ�ӣ� _��qN��Dm�g�+�^p�aA��T(�3�">-�d+�����Ռ�.I4��l-��B��lڑ|ֽk������K����7XYF�>���Ӡ��ºr..��*���Vi��	*��[��8�)1\l5��]��+w8W6�\�$��������l��e]�z��l)j��f�̙]�[K��!�����^�v�S�΢�tϢN�EC�
�;��-f!sܑA������>_	�jۚbX��eH�D�����fJ�r��`�7,�! E�4��y0n��B����LS�U��@CA�4�OD�*��w��)�)QX~�U���Z�J)SH��
�k�`����D�o
�[T�R����fQD���)c;�{0��Z'u���KTXY^	8n�Tr�����Do$4اpƺ��m�/����I"�]?���պ<��DD�R0�Kz5a����Z�.�`@�'��T.-�{RX[�ϗr=l
�xm9���,��.��}9K�rX[�z�Ns^���j��8A�YaЙ_{~h��t��Vȓ%/��dDdS��ټ��}���I2Ԝc���������sj �"��|��YmV[��5ގ�Ȝ������D��٪ä����>��B8UY^pC��14����ϗ��E��H��_�Q����m�/|=���tG��&���B2�FZ�s^�9�X�@���	^h�u���{�a�g %k2�+5��T�7��%>�B��XQT������<.9����โ1I�b9��"Y��~A��bq��V�}m����i�r������\Ҙh5����ܷR��7d\╅�:�]��������7��hIq�9��l:�=�V�7���8	R�:�����hJ�-�+�oa�L�� � ��^��"���G�S�t�l�M�
��vDn׍�������{z�ȸ�&9ڹ+�{:��2W�`�&v�'�w��}�uԠ2���d̕	q��$�-q�2z�ϹP��Gyzj�7Y�,��8��U�r]X�c=����/v�d�9N�~���W��?��T`�n4��5�)8��a����8�Uw��{I��o^x'"��\�ܙZo`W��Xے��S3v�ş-����t*4�d��#R�m��Z��(K%Q�à5V���� ?D ���s3C��7H�g;�J��{����R5���\Q����
����[^��s�t�������x�8��k��+�x:']�}���������_aU�5hLv�J��ԯ��܀�U={c��y�� ��妮�^t5\�&��l����H�No���@APb��Y��Z�-0��xJN�]�ʐɄ#�O �w�1���|�b9���3���i^M�?�I�5��LE}�ms_���H�1Z���|�*������'�\�k��B�d����c�l��G���|C;�f��m ��!�\{(�=gP���D�5�`Y����V�}�[OI�y)CM2m�TD��n>v�cZ�M���2+v��m!��eÈ�C����a����<��{�aHί-���#^¿5�E�6�� �GԨ�4�H'TU}������[���ݪ�,�����$��5)gB)#�Qwi��t�-��)�Ϝ)*��G�D~h�!F�����4�6��9��7��xM>L����V��F�!b2���qoXI\a���rņ���g-�\v���`��\�?��J�j�ܝmB�J&M�0`nc? e�!�4D�b�e�$�$+��#t�6@(F��N��/���@�aS��^y�H�b��!pTI2�z����	θٳ=%�t�����M�`��j(�r�w�e�;��QC����F� "(!SDc��;o�f�v�v&2�	֗��X���i���5hz%WO�2�O{h���F�#_��i������h�34�χ^5gdHdp���2|:��Ԥ�@|�\��F�<����Ri{��=��4P�c�W$�g:k�y/׏,�+@3k���&���u9(�
���*.dL�.W��6c��&! �|Z3mm��}�+����0��P��/��Kq�"�zUhޤ~AU���ٴ��lt�n}��,��"������ƈ��p��Y(;'|����3��G����0.؂<��[-$_D�cj���(�qn�$����ʩ\�L�aɤ��|e9~�A���H��p`�9)'��,ѬQ��i�
ԁ8�tܠ��fPL�~�PJ�U��bmH�..�q0�B����Ph���u:7�a�e��̼P/SE4�{�o���X
��>>gŋrDA*�"�/�,\�f0&汑X�W�`ܘ��7��\�Y������獟(vU���G���_+�G�mc�5S/ b�0�l��c�L}�a��2�̭�}P~� ��E8��;���4��u��h����W;��[�xtUw �K�����փ�!�E�ۚ��8���J� ��2�g�2��ꌙI��!؁�,����'�E~���兣���`�r]�.��%\!��-[%L5B����:=�A����_B�Ǯ�ԕ�����P��n��1Jj�����*�=n|܏�b�t_���sýF
fd����p(��/H�{"�3����s�,��U��f/n�4h�@J�xo��e�'T���'y��/=~��'���nrF�c|�j�s�y[��J� ��r��c�xs�<0���"�	%hRe[��� �I5���ZB�K�U��}�0���6��4��C8Q��H���E���~���}Pᣝ�̴�C��u����wnK�~|y<����s�Hk��5�a���@x%P����:�jȋ�f�U9E��[����4�h��	�G���Lg�-�y�B�#�`v;,��yGw�ڙj��n�����vݨ�����Q��K�&wc�A�0��ʃl	|�����.���X0H��Msr��[^pL;��1�N�~�]��ޏ�5f<�ީ����I��8aY=�g��V,.�N���Ң�r��Gj�Ccq��0�^(�{���$S>J�䜁��� ����^�z����H�Ô2:�0�65`h\f�48x��K�@(��^�m�R��D��%	��>�LN9~�Q|��xj���D�~�4��e/�:ꪒ�ZJZ��'����b��(���䡁CT]-Ӈ�ey��z&��|�x���D6M���3~G���X�L���Pݻ�����į7�� �����S�ͫڜ�=	����7�bB�sk��~H~�su�%zX�	����Kp�	�����Am^����byz���]1�7o�cbAd�Á�6.��Єa�B����&$��8b/��<���7��8��'�,S�%�� <��VtL%��&w�X��`���8/�6�l��7�q 7̗X�H�9-�Ş����<���A%�?zU��ŠKQԪ��3u>YƝh�m���$�D��W��#���$�G�?��	�rl@�N���d8e�pӹy�ڭ�'BAQn@��M�y������A�AtcC��6[8��H�rs��XA]�Ƹ�����z���)����ߤ�t�@�[[�E(�E5-���C	==�Ҫ	5�V_Σ�+%�����g��z�L�	lM%����m?�R��7B)9m��YJ~���Kt߽���ǹ��o	i��ގP���S��B*b��i�'��J�F<��`vh�ny��8��
W=q�N��^3u�~'�f��i-	���p8\����Ь�[�$̯]壬=Gù�����,�\d�45H��8����	���֕���'�2�~ ��~�����?N"�B��o��f������$�����Ss�h�gmx�u��OƮ��k:�'eL[c�]�$�@cۗi���D��C��˝"���1�k��H��E�1���*[�5�{Y-%vP��w�a5�[p� �b�Q�Ic����A�.����c+���C�O(�<1S�����.ؾ��z�����
�&��1�+������/�b���&ȿU��_�j��C�C�?���.���z�0*z몚<��"�lf璻 !&�|R~�cPZ�1�_ɹ�7�������� DZR���<�Q��/�������`�KP�������L�d�>�PRs����7M#7AӤq&4�Px��\����o��=P��|_�59�Q�iM�
0���� c�&]Q�A� b[��3�U0iu����x#�n���]H��؏y�?��F��OȬhY!قV6gtg�~d� 
��x-B��2�{�hQ!��Ýv�[@#8"��![�y;v:��
ס��n����<d�&p�nMJ��5ޚJ>����[1�쮖�� �s�?	9��>�m��|�b��K1p��(��k��L�q~����o���v����Q���r��,�ފN�����o����7{!��%��g�B�ߥl��re��J$w����x���܌�� ��h:��^m�[{V�q���{v��J���s��������͟��^�ID_D5pR���ʜ�y˳���|P������7��)��k�찛�d��1�S�h���Y�߮B�����6�ѻ(O��%⊇�C������#g��m����F2t��T�f�7�'��|��& &�^ �(��C��Tۧ���ӝp�5U�#�To!h�f��<�-2~`Maf����#?�ٮN�L�'A�c���*	g�n�_���%� +�����sM�9|"$_N�������@\_�����%����vO�9����"X�s�?+ D�E���S�K����dO*/Xж*�σ��%��b��yfʩ�x6�%����(����v��D���94�����U���46�2�Z�)]�Z8h��������l/�A~�����oQ]���x>�#]�����A�
�W���TR�V��?�<?�jpr�΋]�[ٟ�y��;�l"̑���9�EE�~���vM�&��Y��-Q�J~\B�=�)�p ��
]���"���-�>��2L�P�UP����Y��W;�֐j^�n�!�Z��)�gF��/���+pɪL�3�?�>���\'�S>���k܎hpC�l��g!B��1� |t�kg3Oþ�����մ�_T��v	����_�U<���G栦6?��h��"[_�;�?�p9���[#�7zi`O͂��m�|q�9�ޡ�C��A��q�CӦ,�p�܅6n���T���!j�1�3�:���>mg0�.���2K�������^a'��J�F��D���W�{_�H��6�_o�PF{_t]a*��E�q�R�Vq`r�������6�b�'-q��`k&��a37ܺ��.�'��pe�c�c].�y�Y$��7-(�*�Ɂ'�D��:F(Z�����&aHmd_)�� ���@d���vJ#mA�K�(&TY�</�����P�c8CZgI����;�Ț"��I=�d��Q�f�ެ=>=��DV^���t�-���W{�hi�bM�e�°�Mt��.�|�U�[�z�k��P�� ���~D��k�9a����_�q�y�N�3��˹m�	�0gu��8������2�2V�&{�� ������G����7�Qre�j��,���s�3�8��O��	�Lij	���X�{8Yܧ�%\�D��|��J�M���i�W��f2�'���п�z,���Opɿ㶘Ј��+��3h��d�1�0�Cl��