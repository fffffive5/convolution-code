��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L����ʩv�*zi��$��SMZ�+��j��]*bD�+wK	�eJ��-��}�BJ�,�=z�޿�I�:���x��K}]��Ǣ�3XZ�i60�_�;EW�� �	���ü�t���T~X�j����9�@��UB؛_��Xۙ�ng�L�s0a?K���BÙ��q!�rAT��Ե���P��΂f�?��ȩ�4>B����DDOɕ�EEܙ���j��j�T���={��h��s�l�ӡm�8	��Np0���8�')�i�4���m�S90g5B����x�P�&q����b��^�^���Б��73W�Iu��궮�ɪ
S�=���y�w���y��A0ÿ"� �~Ç�'}M �E�T�"Q����I�l�HG�[�ԧ܇3���H�	R���<��������-Zy�a�y�����9ew��k�]�%�����VnY����tt���������w@�<tYw��K� ����^� (y��;��-	��H�F3�� ��g�o�$)3��m���O'� �#��VNL������f%ݛ9�N������Ge���\b0	�����u:�����A��;*��.=�I�E|��{��;�N�a�9��ut(�z$�ump�މ5c= $�j�?a���ɚ�`wZ�V�&A����a��hs�@�k8�ħ�-n�P�?����}t~d�>쓋6V�pd��[x������/j���@Lr�FpK�_��� ���_�@�Jr��0s��|B��I��� C�����5VT�GD�_�]l�R��O���h��1ꝼڬruU^�i�w���v�B[̐��3o�%�4`�	��ȴH�T�8������Ϫ���#?$n��'/nl�Y�c6K(B�����W�sl����i}rEb_�E��o�1�G�rw�0U=ޑP�� ���X>��Iz�3�q�7wIp�����.tv��4~}�(�S�ǀ�0�FB�|_�b��<����.�|�?(����aپ�٣~��%)�j#��E�o�����	�n�;g�n����Ց�z�/�Y৹ˑZ��,Y:�:�U�fD<����L�ZG홴Y�>q�r�W�Л��v�.���?��c[��(:&�Bα��G�(��c=����?��4Re�(U�g5�ܬ�/�⍀�Μb^X�]N�BT�Vt� $6�ӷ����k�PV��]���ȳ#M�t��0W�@>	��/�j������!x�U�.��<T����?n4�7�b́]2w!�Х�*���.1��lNт+N�.��T����Bf�����@>Nkw_��l�bx=�I�/cD��-���9�$�=4X0/�	 ��x+T]8�?���]:��*#&��$�1O��(w1��1��7x:��`
����>¶�+��[,E_H~��Q�U����'Q����0��ӱf��U��ޚ�x@vhO34❿�Ԧ��xyR�v�Lt:k�����F�F���g�U$�~���B1[x�cSd�C9j�!Q�I%����s����a<U���դ�B�ص�/,�T�gM�1F6��������ϐ�����aS\�~(!c���5h@��{�)I��y��|�kEժ�h����Zy�M^C|�T�+G�l����_�>��.�:��(r@���e���[gAK���q�0���f��w�x�+�1Tsy8��"�Zs��3��GKډ�}�;>\l��&�`�Q���:@V��V\�=�@j>�	�O�e��FI���/�G����g�0��B^&v� ��?����&���&�W�f`o�7L�9��}���y5V~���̨$D��	Xǐ��H���T��D[9]ک ז�_+�=/��k��7�����-��%
iG�؊�HZ�=�zģ�+w�ܥ1>Q�(�׺Bl�aX7��I4�OK�q�q8�*��*����>����)��ٝ1򾜏(;a�D�#{��
'�{:Ю!#���- qD���`uW�,Y<�H�l�*cl��+WZ�ܣ� e���	�"i�������|q! ܩ]I�3ά�ukT�k������/�r���+u U���ڑ��"߇�Ȅ�f�~�Q���r�ja魘��Ki��x���䍾� ����pM�b����p���M��6��Y'�ь�0�x�(_>38?�K�&�'1��Y+b٥oa��#�N�G�q]�o���5��}�*C��O�;���Sម} �W�L�9�Q�SP��?� 0Z���a�O��D){e��[�-Uf��#uE��ߟ#_�r �)+�wO��B��<��ߙ��Q_s�^��4p�}�B�ƿ�é���)ݮL�A��>���Z�w�My�A�o�#.�|'Lv`aY�K�	F��Kqe�����|S�Yr���o'Ա}���}+X;�3�a?
�O��W����UG]h]� �ևWBJ��ƊoN��B7�y��|ؐ������=�¦���	PHIH��#t���=��\���o��N��1�����'F��ۼ�/A���H�*4E�}�I�Q�X/'��60?E�=BX�)Kpt����f�dP�6Q�a 슡�5"�<�܏����u�`����2�d��\������fj���剺��#5��8���A;k���ɳ{?_�.�U3JB���/>;�}p�
pÆ�J�
8c
��F�)cWH�==C5������4Ϸ� �kB-Yw!���t߰�\6��~��8���s�`丹f�����+�m	�{�\D��.�R��z�Ҷy��� �M|�RF�����̳������;8,0`r��ٻ=�V��k\��,��/dj&����Ϳ�,Ӊ�֭.���=Z�v���u|^���J�(p]%��J��9*�0�hp>�
N��2��0�3yWU�t����+U!�r�qv��8��������SA_��҄�n�*4��`�6=!A����]ǅ���ia\�̇����"7p"�4�7��E���CqeE����Q���VG��Ǥ�6@׻�Ov�б��xB�|՝Rp4�m��K�	%�p�����c�G_Ѯ���cG28T��w���Ӱ��*$~��É����L!��-���I�a�7�:i��n]ݦ�f���*�?'�($�Y��n�����d>q��3��y5\1�9��5�}O�5� 4���)bޗL����(��d{����x0�`~�2�]Q�Ց���Z�=��52�H���=ڽ�	�2�q C�u�.������f�̤���R[GJ�����7iaA�aSK7_'���S�[^0�E� b�*���V�z����v$�j�:�p�}�1y[:�P�-Z٩�1?j��A�Q�����HZԔ�f������h�ūJ߿��SD��;������l�&E��/�E$����9�q�7uY��ÿ�<�m���~)|da�42l4�&j��z%��5��)��>��Y���;�Av���>Rw�#�ww��ᥜ��p�����(%��)P�C��޾\6��w���OV���RR�&~E�U���_�XJy�����fl�_��ۙث��E?�D��|��3������EK�_�K
VM����
�Շ��T�1��g�� �c�}44�(�{������P"Y��Cw�c�X���y�bpNց-��#�i�lK	&�K��*+8x��I:�t$ 	9�ie=��8n�.@o�T7)��7v8��$���H`~=���E�۶L���P��^)�D�К!��!P�/9�oU���ܴ~\&w�!�2K$�yꨲ��1و�{_ߵ���W\����_5a_qJBv;|c�KC㋫1�)̌���9��6��0��s�m�c����)������L�nN6Jf�4Է�%�&^��Nˡd�L�E�B�o+R��s���X�H9Л�_�X)��ө���@��h$1W@��8���T����ǋ`���6��� '���S�\Ħ7<�s�r9�ZИ��HC�r�B�MX�OMG&9���s�6����I�%�	5r�:QlQ�1P�ٸ��r��a�c�`_YXY@:�=9ׂ��{��f��"����w�ޤ�ُ��N�������V�#��o���=�{���D;"�p�@*����T����9�`�e�fRUЪp�SX�s{2X����L;�t�Ɩl6 �N`��;��v��@���U&��2^�6����f�m��};UQ�.1����ӐM(J�i/mZ������T �g�m��U��4i����>�|5H�{�.?p���=����!E�<"��7=t��kPd����ѻn�}�0y4�@$�̃z���$	�Zۄ�kP@|��i�j�Ҙ\��w�XY�~��
����&��kf��ݲ��@�4x�%Z��_�����E=���yQP�V�''0l����~�r���b{�|h�,ڃY�� xZꆠy]���u����.t؇�<:�!X��-,n$�PM<bF�CgT%�y�ȓI꨸�l@Y T���<��W�DR=��ʠf�k�ŉ��M:<f�W��$�� ��<�ϱo���H��0+�?�]ܨ��0���0>�nS*�]��3��f4{��Ǎ���{jXU���hR��EdNt'	�_%?�o���0��k�����~��ѳ�Z�S�9Z��Z.n����l����#��Y��3*���0^/�iN��ؔ^I�>W�p���xJ��k��j���dx���#�r���AVNĥ�X��v�R��m6��+�1�|�{�H��H�ӯC~��8������D�����1���R�{�rpp�m!#��ӹ�K _q�_�_-�0���5�aÿ���K�oTU�'p ��\���ߢ;o����!��O�'���^'�|UF���?J���e���e��3r�Or���֌�
`j��~��R��!{�)�25*y��}�����r�d��:�v�\��K�D)�<h�xo��Ǆ���_������4��O(w�mD�C\NaE��P#��=H����s� Mqg���h����1�b���+�Q9jr�����zr]�R%�d��hO`�"�v��=�h!�{�yB�*����<�8q�y�$
VO	�l(�R�����
*��]�W�E���=� ���n)7L,���#�S]^��A��'2���ꐜ'�aF���F);(J���.Z�V�@�aDW.�W�b0�>�"�"�λ��W]F���x�<�`���?��m\��v�3v��+�@5^�+�]�R]b�]V���&�!"l�/2��(ҿg�]���uы�g|7���?����� ���;Q�@A�f���%�(�d<�0���*�r����1M'{ZeK���9C��f%l���P��^�ё�w¢��ޭ�����[�����JU3+��X��UN(��3�T#�i1��%�z����f��hYqװ�B�`#-�y[�"����	��!��9���Q���:�F��2$��<�w�
g� �0�i-�/1���$9a�u���2� *�=�C`J�!0n��X�4O8���aU�����$��H��Pm����[M���^U�I���md��GP%=�5d�.l��M3I)5�k��-Y݄RU���
S&.h@)%�SG��W^��ls���(�YP��,�9���q�։%�ܓ.����Q����ד[H�Ǚ���H2�~<��>�$f�4�gz��q܁��k�j;o������>]W� P����Ec2�GC���yhn�@���;�g�-�ϝ�7�/olW�V�u�ⅆ=7|q2�G ҙ��"��B Y���vW
�K�,Q����jF�a�zGX��b��p��g?�@�������-d�	�#�a�k��(h�#�0�8�{ppcû.ӧb��koJW�.�)���c�e�W��Q�IEKj�*)�R��6��"�-�޴���5V�x����B�����'�O
�d=��g���olM��ʙ]=o�(�th7��}�1l^���/����f �(�
�>!'��9��>|�� �h��S�ba�P�3S�<)hL-��*��j-�Ĺ��⪝�����M��w���m�b��$hry�h�n�J�U�؃ ��1���_�B
"�ZY��y�uЗ9g�l��|8�������(,�PR1ҚWĦ���9or%��)�0����{z\ö.'N8���u�p�[�K�5򛃫�>�"*����c�Sc��r�R�eH �������<<�ɟ ����?�psF	Sh���y:�J�ˊ�=p��tG�b s���ߧ��͒O%_o1+u�	����u��?��]K����X��SY3�V�-����nx"�,�-�7�4P���*�d���b*���_����)�-�J�I����/�j0<a�VfWԅ��o�xNXs�N���)<9��a#x�"ΦE�mï�G���۬�r��b�c-)ɼŜ�:�3���U��husYN4���fM��F}�V(�K8���ͼkF�ۊ�΁�#�t�x	J����݇d������l�~�X�O��Z%��X0�dCsR�[l��Ţ���u=τE�R~w�$����΢,�����O��Kwcb�0��I�tlz��=p�5�����+B�u9��`���>�*���~��}Ls�E��i=�Ȣ� 

��0�95?��qqԁ�k�P�t�`
�a�B�%6��-r�_[� ��<d��w��f�U+h���ۏk�[�$'gͼ�iWf����P� ԝE;�na���oՑ�wwҌ6�+A./-��{� ���Z��g��e�Qՙ�L�<2Vk��4��t7E^Ժ�@��`Vp�"���;{$��rUwd��s9{tL�}L#��J���޹X��CjC�y|���c�,�K�a4����1&�ۥu �h[�2���t�ݛ0��t3�r��.�g�-澖X�_bϤ�Z����[�6G����~�Vet�:'�׮	;�=woO�di��:i���!g ~`���A�W6�W�k;�D�
v{�֪��U@}4v�!�K�8G����V�^�L$��
kiF$a
S�xS�̸�N*K�A�3��]	��b��%'�wCY�&eW�+�J��D�c�6$j���C���_���B'z���ۖ,��e|�������i�^+P�iB�����Ep��>��鞅���}�>�0sb���������88�C�}�y�k�W��Tx�U���4.�j��M��C�S�@@ߘ�3�j�ˡ �^���{��^��LOPB�O�X0���N�o�+.����c�Q2��{="nL�[Z.�F]<�Q�-��.d�R3Ѡ�����զ�yQ�x�p�e�ǰ6l>�}:5���L��.n�2T�����Y�h���_�r�U��t�Ho�	q�?%5fd�$�cHH��L�щ`כ�^�u�q|�و��U*��G@�(1���_^(8�S[��gԽ	�P2�|5��=핋��饴Z7nh��N�ٗ�ڄ����������z �l��3YP�L�;m�]�`�n�n���Q��RP���N%�c�n����̥<������b�[�j�ɴd��)y�\�fh$�qr��p{�|�p�L~u^���i���Hyv��S���f��3������q�J�gE�t��O��u˂l �	m�-�c:p7��mc�����M�����'�~+�P�S,yb�S�ѵ�L:�l3v�4�x�_�#���nEg;��G�cI��i=�� ���0�|������L�T*���]���r%\�������(�l|����í�������N���J�y�8�%s0��#Cw��ES\�41ɶ��R_���P��&a@?�b�\"Q�EC����-mܟ��!�*s�[��.LG9�ɷ�^�Λ��������=�,�A"��p=���҇fށ��9�!�¬��9��W�b?S>�k�ǰ�>%�ɰ��@;�h�;�wX�"x�v.b߹�FXm |JF��@�3���Q���P��`b�R2O��y����f�A�'5��0	�2ҍ�.�P�֬C�]�GŞ�������:t�r��	� I�;�k���>�q������3���gv�/��g�Jd�ʆ���a�z0�º�=����c�2�#W� ��]!WV/�QKICN�O$g���y����܆53E+d����3;�4��	��g? �3 �r�k����:��N.�b�P��s��]Y�U�ܰ8*�X�6ަ�0X��0�V��F�6�p���bQ���=�އ���GǄ�k-��`����MU� ��&�7�<��9�a���f��K�u���$�}͛4+6��{"��y�|�C��KP���,:�?�l��V#WX�-��[E��u�3��0��E`�vF��|����P[���,���&�:T]��e-WW˼�w�������E���
K����������Bx���G�H��A�5�ԣ[X�!i��my�{Q]B�u4Yj��ݐC�mL9fD����h�H�:+s��b��f�4��y���],ׄ*�d2��jP����R"������|�fciRHA������EN`v�X'҅�*��U����Y.�]�)�\�/J����g��k�Z���}��(��h��N���{�3Y�L��[���s�1RUtA�dd�jDGJ|����)�(��@Z��}�#}���٭�׵�Mz�
��"����'CH�<�ǉD؏_?eI����7�B>g�}���=0)�k�蹥��ȶ�����%h[���̈́z�bxL�bK���N�(2g��U�F�O��%:>�.�T��K2��?����nK�~�q
Ht���C��� ��%��
��E�&��ߣݕ�-�x8Ek�"���R��p�R����K�j_�"Oo�v�����NԳ'Vy4���z.},X��uِ{����oe�ƙ�1� ���g;�,
��A5`���K_c�5H����g�ރ%�N)��<���덢n��c�h�?��$���p��1�7)�$���H��h�N,��$ i���E��CH�?��I$� }��a#�	Jp� �8��8���',�id��h�����P�GO���@��B�!��.Ky���%-�P(��%'�z��O��^�����;Ձl�OQ�0�: *[�"����P�@jK�ԯ� l��Vq��1���1?�QH2���pt-���X�˕�GxN�s3)�t��V������Âr]xGz���CX�ɭ�NE�I%��>�L���r���Wd�����N~?*7|��ה��e>�R^xM��K�&e3�� K�`�Xz�����;P�-��[7&J�>�#�A��r�c�{P�Kp�@�@j/�����"��L'�@�#l��K��s��~�����{]�1�,�?ܐ^�Kl���\or:8 �����=
Tg��V���	�R^R̽��Oc��tA~�!��qB�輦�� �(����>�|a�4b�l����b�r���s%T������:�AM�ƽ�@{������� %�LN4|���TᏍ�I�/䶬��Z�ѸL��G���ņ:���'��o�5����ZS[-W?����'�H��Ry��f�A��B��X���l�Q�Kv�uS���@�	H1��r�M姧<u�MdE�djU�Yj#��V���T�d��������:v�X��TIe���.�F�K��ı3�)ވ�xZ�4>r<��gZ����3<\����;�z�8&�������u�V�n��ҴO'%J����s�𖚄O�\F��0!����nq�_}�ŕ.�pd��1i��z�H]y]V�_����2�=ڴ�e�
�A�F�"�M�Ki�b������7�)��'��~(�X;~�.�Z8P�p�3����v+�j[�d)�8	�P�������II /2��ۙA]pq��*�&:�,Y�'߅μ-h��CU8]~��N,ID����e$�?��ܾ��YHV�5v�fp�%ߣ.bo���*;H�k�=-IU:,��d���>�#�F�3��?t�]�um�5�A�+G��G�[]�\�-jpUZi�tž�R'�N�z�Ad�H��d�	&T:ο6�{t�r���$���u(��*>^�B�R#e����#EE{�^W�)���O�sO�m��^JA��Tp�%ʗ�4�*W��u������Ԍ��	�kS������gh[
���C ֎�V0t�70'�5(Tm;Ke����V�ap�����a��M����y�3�6����Iq\%&7ލYXqq4�r|$�l<>��XA�cKɳ�W��U��JG?R��-���Y����<+:�j���v#/��#��^Ab�������D$��|����h��n�d�U��?|��s	��T3�L���D{6_($�f�ڸ1�h#��3)��VY{�ϟ����/���吵���c��&1 ��V���Bp�בGSS
������-]G���K�`�-�g�]Au{f����SK�;����3���h �(7 0z�ji���?�	p��߳�������GSX��/A�1�r�n�[�c]�Ы0������7ț� �#'��h u���lK�����ܿ���� )ͷ�/�wyl�Z�f���d��E��?.M�BR���Y�n�w#"���N�lyh��zD�W��gTx�����縷����C��Des��s�-1�y���|\@/2YB6PX��5=�� sF���.NLX��@�b�ŐBL���&!�$�3��̤t��U�M��K$��V�]
8:v4`�f�4#$/6�E���tN4D[#�=��i�H��X\���������w���u�����{eR\�7�mO@�m1aI�[��A�'#���������dz0:l����;��"�#nb��lg,s�6����A���jvb�h�d�}���* ~�.��Fz�ʸ"7T[���.(%;O|E�i�^��eܮ��U`dm��H)� !(-���ՐcC�IX6B��mq0�7N��a"�r���[`I�²S�N�2{�3Qi��V��̊%B17�W�Շ���97�ꥹk�:2h��V�(��]�%g��5�m�-��
a�g�Q�A	�D�/�!��]�(�V[,t��5 ��yQ�֘4�2����sO�&8S��(u�D7���н�����!�EJ�i���7}�P�m�^�p l~�ߐ�H�du�A4f_�g�|��ڴ��7kW,m��W%΅�
�~�h>�}e՚�,ރK��j�Y�d�X���]aM-(,ty��v���>�T�c(�Ԃ�?<�{����I��:ٰy���y����8rف�>҄sU5���?��w���b���BO@�ӟ���B�s�-�@����=���Nn��,�[�0@�H_�w���ӭ�~M��Bk�̃ă�`�Bc7Gd,�<n7�ܪ�]��J��� �!�J�0��ĩ��Ы���R?g��W�u��_"c�YD�� ��]�)�]2��UsW������1��I�6�U�]6��� E��TjZ�j8�� {q
�S׍o��N��p4�`��O%������R)�i�� *� �#��)���y�(�n��g��i�Y��nq�c�G/��q�c��S�G̯^YN�N-R�$�}�Q��?��5�*�p"�<�\*�����\�01�As��?�2�F��v+����Ĉ#�D�� ��Sc��KS͗}��*P�i��b�Oܸ'��+����h�-�3(���Z* Ry��aH�2}�(�)���݉k���SA�@�E�����8��Un%l2j�2�I$�k�2B:0��?�Q�\��wd
�݉7�腝�S����ѽ�����^�"lWZ��\,�$S�!�EC�l�)b�GEh��|b�~?^������5�>Z!�6@�.�Dqڝ��g��*��7���,Vw�k�fv�f�+��v�͎��`*5@���Ycn�9����}�0�y�ݶÊ��u�8��d�'�Ͷ!Q%0��hUgT���^$UN�\�E����
Z��䮈�~]����d�ׁu�r��5���ao�q�d��G|�Ι��0̲�&(d%����h|��z�h���z���]�u.c�q�O���MS����� {4B<-�8�a�������euԳc����f�{\�t�Z��tG3��T��>5f�c�T }j5'Ɋܕ�229����P����p9�_�L<y,���e/���`��ڂ՜*@.���I�=3J��=�'�.��5zlI���C)�h��|��KU��8��s~�h�+P��7��_b��ie��-��GCb��3p  [ZC��t@�^�O�O�N�K�����k�Z���s8�Ow�9<�?qM;V徧Em;�b���TR�R�̛\�L�Lњ?(t���XG�%eI�z7JI*����x�;d$[!��]��p�k0��uR��,�	*J�Y��nl�Hde�>S2�~�Ǆ� #B'�[�k:ݔ��� P�^+���L|ˌp�5c�A�}����%';�ѷ慰�������e��O~���>�~�@6~���{��M�M�c
S}I�wU��U".�:�{ԑ=��Ė���4q���2��#��J�;�I�9�R:�Du�i>Gy���yd7ܥM���r� R�?�J,:��Z���|%H���6���E-�)E�a�*"�4�J*�W-�n�}��8'���:�.V�� ��O���/�i�3���̒�SJ�ş6��A��Jl��|�&M(���	��T�Z��#95cm6�R�+,���?�=p�A�3Ս������Di��E3��߀4�� ~��sX�V��Իa�bjȐ�scq��2ue?��2���!���D��Z'\}=�I=�g����:B�Zǂ:J���5'�J�F�!��r� ���~g��~�I���Х����MԅC���P�"4�8����e�X��+�����dp��H�ya(�ԕ�A'�dqy��:�hUW�,m����|����e�$���Ng
l�l!��s��槎d��Z/=�qH��K�3�ͳ�R��J��r`2|�gyݞ�n�y�K��`���iF\��	��	޼ŝ�@9�/�P��p��Z+�\o1"T�����!*g�?��e$���i�y(���u!J�Eo���X��@�O�~���t�5t�M�&�>��ӻh�a�~ߣ�C���nI����-�9�zLɭN ���L��Gw��$g��YS�f���W��%g-�h�\.M)�zyb2zp�&�����E�� ����ZQ�K�Z�9y֥A�\ާ�Jf\b�R*���|�4rf8�����2� �Q��|"f �<K�� MI���7s'2�,��c�h�1Y6�g��<�����UQWa�K��n��`Mr���"�� �G��E�N�H4ߦ]^����W��3����x|�D-!��%˯�RM� �Q��^������}N���e>ʧ"��:�̩bE`����Ρ�|9󀠺����Mt�����1����QV�J����Q�N�D)Cg�����M����|����?,/�Z~.���!�h�PWw��V�V��J����8�p�	1P����U X�>���#ɍ�v��Q��w`Ok?V�V����wV�Η��{B���\�b���*{O>�v���q�xvDtޞM���������t�.�\� ����1��Y8=�&�4�"��t�o�go�.͟&�.
ЩZUW�Eץ�6dh�uǒ�AM)_��$,���L��lS�,&�R�Iu��~�����@�B���u�-�^��d��f'K��^�^kb�h�oޥ�Ȑ���&(;Eߪ��֥
��\��n�{ y�I�9����±��B[��|pƱzۿ?�G�cm\�^���\Z�������������HСHY�a-?R�h��Z���MIZ	�����h3�K��q9r��:���3S{,,�����(���2�ǔJ�*�����JYH[Z��J�f2ipgSg���7�d��J�nЯA��Ԩj�2X��S����C	.��YL�b�GW���v
���`E&���W���Č<ɗ�§L���M�Z�N=�� ��b���t��Wb7�gۣ��3~���Z2]Y���,�T:��v���}
�B�|�X�`���Jɩ]a��'W�P6���'�(f��g��s[�YѼ}'�^���UD�Bo�խ3`�Ln%�&�M���\_�)��bM��2�>Ũ ,��(.J%�_�P�N����:F>��Q�!��yz���_�I�ښ�A�.2G׿|Dc{b$�4@�U��k~ad%�Kͬ7�:R�:��(����{L>|��������{�
�>�\*/�]�{�o�⡃SY/T�l��i����G�M���.[S����F7b�<-F�[�x��ʏ��˂rH��g&���yp��1�{�o�B��#3Ȍ�K}�[�	����ƴ�\�2��q�
[\�c=�S�+�0QH��X�W^���f�L�Ǩ�l�I�|����9�mɹvҨ�����w����9}<�ƍQ��<s2ߩ��.��e��6rk3�N/ E�:�T�hČ��!"%ƕn��j)`�9QU�����f�Cŗ�]�K�O��1#y@V� �I�C#xXD�2��Ϝ M,��ϝPN��
�rŮ7b���4ү�9�]���p�Aa�L��61�\�Q �АBv���n��N�	>���j1wQů�U��(q3q���^B����f�_Y�H�^�,KdUT@��89ճϾ��jI֧��x����%�K���"{���-�t�_�8Uz�&��B�7OKN��Qȹ�NK&�^V��1éFG���N�l����	X������\>85�t�_Ər�� Gf��`l��OV�]'{��Z�i+�u����8�(�>�ªVG�x1�(0m����.� :��ߎ�Z�^5�}J{!��f��,�!y��s�41�[�S}1rv���6pmK�u�sq =�3=7�p���%a��q��it܏#]W����f�d��|�h@xY�?Q<N���6��r����-̓�!��7�*���Ȅ��(��]���pa0��S��Ӕ�h�J�S���hꢦs}C��E4��7�L ���|�����NS2���t�F�2��|��q�-�g?B;�N���� �F�	�����+�<��m��*!yP�#�j&E�܉��GZ�̺������78KZ��@�S ���{�~��jb-�� �k�Y�}���.��P�JR!@���۝�_:���e���������C����nb5ǆU����mᬲ��.`��^vl���%2W�}��� � �v�a�+�Ϡ�A�N�V:����Ш����$�ڗ�a�d��$�(�ܶ�2�-�Kl9xI���Ȱ:RV{�5��Y� �С՘��%N���0��UǾ������RSj��M%"���O�L/���~�F�>f��KC�.�ފ�~���(7<(��f��D<x�Cka�]�泅�J�}���z�ȚE�̙��#U�mr����\� ���&��M֑���eɶ��y�ި��2Tbs�'�MK@��~�C�%�Ni<%¤)����jq��<��7������&�B@x�_�X��$�UA�|
p�
��ї�6S�@w�zzƑ��^�1���j�qLRI�T���\Fl�nb�x:eDL9w�F����q$��dL��	L�,���T[l.�<�t��&���c���Z�Ʀ��P,K�:&,V�&n�p�$|��	%�V�#;Ջ4. .̒�Mc� 	�6�E<�}��biq��,�w6�N.&ӈ�k��p�*hA�����s�=�x��uA�#0*�ӏ�%>A>�@16�fr9��I�
=�[3f��Uz��2	��E�� H˖�j���>!��&l��ea��b��(р��ҩ���|�-Q� ����<������� ���j�����˘�>U�2~�q�j�d�J�ȫ>:��}r?��|���wء$����g��HY4�8���拡w�Q�j�5Ȗ��=��도�wZ�l )筧#H�غ����2bJ���$�a4�`qR���.��ޅ@�ҹ6�q`&���-9�[+��>%�8�3�"��H������3��5a8���Z����f��V�ʫ��|�^�a'~� ���y�)UV�o�����4����z�E���J�p�j�_�5� ����e6�c�y��س��%�c�D�/����yI���ަEO��A2�-�e�/��"�_b�f/%�x��L����[�9W�ޞV������q�-�)繼�k~l{�I��sP�]	]�!����ֽ3�|�X��^�8�-������܍s��xd�V��4Wu�L��V/����/�>�'�W
O�B��[�h���\������Ln+�����W�p�چR	h��&��CZ�O�rꑻ(U����O����'��5�M��t0�7Y��s��*����͵Q9\���%��c ������Qn;���ϧD�e��)���N�Hd������s�"�<�%
�0�c��|#rH+c런��j��w�FM>N�H�ߧ?ɫ�{�Q2��B�y"���U���fb��{6���A���_�~D��j���)���i:�}���pO(�3�^�>��me)p�p���S������uŴ`��ӗX�57���Y"��������"�n|.d4��*}�"S"`'���5��S�P����;���*�f�г���W��I�����$wA|h6�RnkVf6�q�	��J�Ӯ�\A�Q��jP���\�!>��;�do����ek{�S��	w����s	��d��q�y��n,y!b2�e���8@"�7� Dp��Ia�$M�߫W�U�Ϊ,A���};�9���rWr�t���F�(,��J�����G[��5֢��ADhMU���C�6Q/$E|(c0����Q+�0�z�J=��k��n@XSt���Uw[�NB���[�+G���]�h/�%�iE��(L�����B���b��f�����Ԃ ���Գ���G�����F�u=�,�o ��Y���5I�t������6Z�#h��3��=w�҂Q�1 eR5�fֻI�"銁'���7����c�r�#��+8>�3�� ��2V|�"������`}�j�	���eʊ�'"ꌹ����Õ�?q�*����Z7�ǵSM�ܟ�e��j\@vЯ�J���0�a���3�,o�z׫���mz<*!2��f�<E
	���D9���Ǐ᤼�$������ݥ�P0�]Ē"ݼ �L�BHE1����P砕<V5ǤZ��e���VDF����X��J�̙
�UQ�a�58]�&⽷-�=�#��.S�ݞ4X{�]x�"�8�u��0lC���3_em�kcd�v0�1| �[�!�"?0�:~�Ȩ������az3�E��<K���Lw��\��	u'������v�;L��A���|���MAL�&��)����ھ�,p]7z�L{�|��z��	�2�Q�B��-��N��$�\�kb�!�aB�ϑ�߻��]��{��&�3�|y�.��J�1���jz���Tj}����g-��"%��\�ݏ����nB���j��Bš�]q,@a�9'\��A�U�_���{���w��t�@��BZ�j[~Q6.6
+��H��d���U�<P|��G��J��0��&�W���wcJEp��9�ڬ�<������Cu�#[�(ﳷ�j��}���fà=��¦%{�����9����fd2�p�-ǯ�0t�N���6I���9�D��6�Sr�C@�;j��{��y!���-�3���A�����
t0�~�W���B��z�u%�,��Hޑ�7���(Fd�!޺w��d%���C[��*��#�ey�CU����ZxW�lu����(����J�A�O︊�kոN*Jm;�c���=d�s}t_2�?򥷅� �>�����'�v�S�,F��y�����o�s.V���ϙ$޸�ړ�
�6������:�5��a���
�T�"�3�Q�r��O<���9��l	�2�t���fX��-6j��G����Y��SZ�$%�Wm���8��Ԣ��@�Кn
�TȾa?Hc��T(������'<h��xK���W�P)�jp��A.Qms�Eٍ%�_�/]B��f4P p����/��1�=�O��ui�&�ѿY(�)�:���/��;C�Y��ͬۮy��a���r�Kp_�!�p�U��Q�A;7pwT��Q��D��#�m�h��k�
��~�N�4��@Bh3�{g`GfF)��.�p�aPS|��@i�ʏ�m���J��}{�o��t��*�`��=m�snz��}k��(�C���s�g�m�s �6]�i���@�E����DRn!6��_��� �X��t���@�x$���.ґ�R�e�̣*EA��](t�'�R�	���Ż�� ��Qµ�Jl�V:��o�%|G*b�V�vo��$(��xa]b{��
툠�y�����0�IU������ĝa}W$�'j�R ��\ {�r;��_���F.L=l�U�$�A���&�Da{�*/�5��2�U��w�fy/R��(:'���V�3_���P�h�ݖ��|�jw����19���c��<�i��YU4pjR�5��O粈`q��s,�l3��64�Ф�:T�xW����)�����r;z#'��S�6�Q�Mb��� �����¨B��P�W�]�����M����<t��,�ܾr过�+�ݩLۻ��%2�h�+LK��'�5����a��fSK���g[�&���oo_P����Q��P>�	��7���]��(�~����n��Ū[C<?��u�6���:�	����ָu|��&y7�F8y#�p^77Y���2������I��>�� ����?̧	�یb3RJ}��Yt��L�#��X%Js��G25�WL�!v��#��4���.���O��O���"p��r_-��=]1tV��_�P&�En#�P�$5A�4~�����I���Vq���yT��Xy�ٰώ�?t̨hm��OZ
��Oƿ����	?"��I^�7�yi�#�U�S�	NE� �(�L�2���� �����y�\fD�|� �v��d=�:������i=�%���V��*��*�*��"��g5r7��G�L=0�ǌ�@@��*��;z�4�o�f�:��	�&�Ax���<Dn&%n�`���3W���&Y^s��U������Oj�^�����MD�H�o��s4�~"y ��Y�0{@<:G��ħ'����vv~��Ԁz
�R��Q[�j�����t".Tr�_��p�!��U�7�+ڢ�+c��>:���p�5����� �C͑�Z*9[��6�m*ྉ4���"Ʉz90�Ɔ
�� ��c�Sτ0G!p3����&��\�����>��;�?,^�c>Š>B@�H&����\n�K'F��밷��fA �B��ܲ�!�[w*�4���#��� ������ H�ԟ�/@"��0r�!�v�ͅ��'�l�]������nx��WO�b�(��ޅBB��{�W��깷} ^�<�Y��lQ�W�h����L�\e��
=��h֐gG�<h�Ƽ��N���`ص��6Q�9�73BB� ��)�%�3n!�m���"&Bl�����ڽ����Ʋ�s�����Ka���>ƅ�<���_��'?�ؚ � ��٘�F�eOXg��-Y�B���n��|��V9[�-04izO$��
H�J�8����H�c�J��.K>��e�i����v�Q6����[�R���w����z4��x�}�-@}����0DO��T�g���:�p2]���nת׀�R>!xK��Xݲ�ts�	$��Nk�kEX���UA�&"��=������*l���]:�r�_(��x�U� �V5���#�CyY�6�a���;�*����"�;UH���i���9f��a��Ws�QD
i��2�i�y˭��=�#��9��;�/0�ޒ^hnY7Z�-'!����ƙj4��G�oK�D��D5;�s#]��L)�M�W��i���y.���͛ٲ���ԙ����{z���w$��zoK%F6.�Wr�Q8ґ'�Z��m|C��@���E��8������o�ou:#�_��}chՁ��d��+@ͽ�07�<�cI/%��1)`$�1�1cu���BzE�ɴEeYQ|C�F�a���)6��Ѱ�gG*�q�XԄx1�a"�n�N�wq�OMV���[�G� 5%���
+���.�:~��rZ�����t}Ia$O����LG8=�3s�F@ᡰ#ViI9��c��ZVYdG�,���K�Z��Rn�?�L�AB��K�����CȻW���8�MP�|K�|
�!O3h��rY���
5�+�������2�uG1�?OC�D�M�tZ��\#a�:���o�a��N�>��56e��bi*�=��@Eْ���he�S ��9�8c�X��Ê�V%s?����j�s�(?�ɡks�ُ���'ˁ���K�/��j��f�����&��7HB� �GU#�C�m���+����E������֤�֭V��ىq�oJ�S�d�9�g9!Xh��'�鸸u�y��i�̎�=��Z�x�/�Ϙ>��[X6x��BR'T�a�.��@d���W?��5�l�}�.��Tyks�5ǅ*���|�P��:}_�Ť�Pt�7�iT�xB��Y@p�aj���eg�rL�ɪ���|�v���~���eOU�KW�>��I�����m���Xȥ-f�C��U�X�Hq���f3�<I�}F&xi�|1��8ԽxK��N�����Q9��{m�U����~,�ǚ�3� � ����ۭc��U��y��1w
#Ke��B ]��E^_%{TA��� < ���㌨��-�n���.�TI<(��4H�7����
�u����r�$��QX�B�_��՘n���f�ٖ��t1�VcԵȴG��B����y�1[��*Kt�1��8���_����W�r�fY�Uʼ_��h�rP��b@�3���!�.9�U܈�E��<(p���tbV�K�O�i����Ry$�#^�>�M���-�D�S�@ޡ����A8)�r��,:1�|��)(|���Yx��C���1Z�р�	"rX�¿<��ʁP	��D;I-A_A�C��2���ϔ�4��CX�������tɏ�W����4A� pzY^��|�l�%~̓y���A�Q�|?�SF^������IS�z_Ǽ�L�3��V��?},6w���߻wŀ@~_��7y�e7R�����NWZy�3T&/o��b��:�bl|U"L-��w�E���9����:Wp`=/G;�β��=K:�Y����������gZoJۨn4���Lo���hح�1[Rm:��B��11��������,�ҁ���%��t�$�/_8���@�(�9����[�'�t������������t-�N6 ��C��#���0kD��2���a�gZ�3��bs"�I��7�L+]$�a����&����� �3;˅�Bh���E�`4*f�����du�F	���ތ��8�':�Xb2��J+*�5�P�iW_����e�9\�v�44��@���%b��j�ܣ���Ԝw8�#�M�D|�Vp/����`З%�N�-�wlc�Y���6��`��u�>�}š�JvגK~9���٬x��Uc��5�FS�8̸���}��1z/����;�
����A�Ěm�m+#�I�/�X�;1tZ�K�.c3��)�96�����nKGϖ.U �.��hPި��7��D8 w���t��=�i�����^��,G�H4���7�(M^��"&K�hc(Q3̀P/Z/$���^E-�R�5^��{N#�v������7y��V���M2dY�tĤ��1���Ylj�dm���n�b��.�[-v�v�ia�[��a9GT>�j�u7}���HQ�61ļ�N��6��+��N�>�Q�V�>�D!���1+ 1�8\��8��W<����}���=�ذ�~�k�n�H8�27��ˇh�vE6�0��Iɂ�H���ͪ	rS�¥M�W��A����P���W�?��Z�թMz�~�S�Z��/��ӕK?��ML���A��T��w�G0̉5ሜ2�娭�߿�@nۡ�������1ʒ����gs�����DvY��ќ�17����kj���1Z��o�h<^�������g)k����������.����,1�������{�|T�y�z����Bn�P�^<�V8+)�J����ŉ�5%yr�;~&B��-4�8�%����I5~�G[����9k���r�_�fQ/�4�������CT�X��n��T�5ېqbcC Xʙֈד9�`�	qH�0|�{�)������~O�jF�����Ը;�IkaѷS�{_*@?��,��-Xk��d,�� �\FI�#���6��ݏ��[��	FП����oF��@].�D���7�!h(�ܢ��c�#�	fպ�����d�H�zWl_�������B���`�cvq���̘v=R4�@߃��28����-	->��L�c3��%>c�h(�Ou�Z��W�5��ڇ�}�l54���\� k�h&"{
-.d���
u�z���8�`q,H�"��&c�P@�z��'�/G8�"��lԴ�����3D���آ�5������u/�n {r�Ш���"5g$����N$�S�<f���G5�b�����G���^[��q��(j�@Ʌ�q��7�X�id�Bnݻ�� �P��`�ё���4�e����˝g�(H�����딯tβQ�'a"*��B�+�b�:6H -�;���������* pb��z*i�C��PN]�W�,;���|�����2(U�2���p�;��7a�Ѳ�MS=éU�A2��OwwfG� ����}��7����:�ŏg�kߏ 'I+X���x/u�{��5>����m�3����n�Z��i�O�gpF�]-gܼA��e�T�<�iKVw��"y�?g;�1o��$�I�a�����v�4 :i-<�ӁMf�3rg+��n$oT|C�F�!Nbq��spE^r}˫2N��^��%�CYl�˩	|v�+��L�e&}6����* "��Ӎ�W�ۦ�鎏kW�49G`��n�5�s��J����P��>D� ��b�c�*Q<AX��c�?:�/�&X6���0�M�Z�������T˞�<;�E�d��|Q�d8�~�����W�r��I����&���v#<�T=�)�΋~I	u>��(VRN�X!�aE��$�&�lՋ<�Uv�R1D��̮%�C[�ڃBa70��F8ZU��{�}���r�Zf�׽�5�䒱|���*�X���sp ep�7��f��Z��`"e����X�n��Hg�������\�p>��5�N���R�� /D|9�Ǉ�k�~)}���7��z��$j�4kܬ�i�J�:�Q�Ԭ��|��4�w�a	�E�sa��E,����v�gX�^��K�m�E0:cf��n��v2{�W�<[n2_;d)0�l����b�E�3e�y�!���Q$>j�v��z����:��̽�z�({	����~��C�ar(��Zh���'��u��T��I�֢f���BZ�(��覑1���&����X%W�v���*�쇝O!����|��p% ��aߍ*�E�ȻZ>Z�o�vp@���.c,+���q
�&rҝ�^��Nˎ�a�OMih�Ā�RE���:��C��"�������T;*F��|��r� 6>־ �/�)��,Ixe����t�#<g�jVs|f*��D��~A%v�#$�-S��ﮙ[-_^�(��@/��K�K��xX2�j�S�NGs�-@�9�˩�ʔ�2~���}\��v��1��)ܪ�W<԰<�˘_�m���) �ﯓN'��5�������}@��$�]=�z���m�W�i<{�X�����&!D%R��e%�?k�m�I������Ԇ�]���$�"�/���d�6�'�M��!�������O�bν�?�Y�.My����|["�0G��0�2;v�N½DfXrP�3��v;|/�}����J��R��M0\�zbQ��T���g2����NԪz��`��t��s�y�K|���%�d�:j!A3���U����R*> =���[)��8	���&t�����uݟ��V.��p��V]k��$5�FB�23�J�@���mM9s����O���q��"E=6!�!=Ԋ3咧���2)t4'|�g��_�h��FU6S�~�?v�|s��2����o�b���eF�}]ڞ���/o�s�=��l�~:eE��EUf�>W��
��ɠ���ǆP�b�ÆڊSF�[ '�S�E+�3N2�]o�r>e�5Q��*�I�ݢ�f�����'!AڐR��'�*s�1�[E���̳t��^��֗�<?��oX�����W�w\Y��.]n�n�2ip�M���5jT���d��i3Hj,�sB�O��~D[D2����A�Ch�{鑏�f�`������� �3Pg��V;52��4��P_�濨Jr�"fF��D��!8zb��ʅk�{a{��Ղ�yB��;�H�YV=��ߩA�:sy���)u?�
���y`$ӟ���VM4q�03�`S.��t9��st�o3{�k���Sk����^ '�q�_�S��է�C�<ց���>�Ѝ�$�R��C�Щd�~|��=�cE����(�![44���&��U��wA��ή�n:
K�~ْA�@ؐ�<���ثR�:���񚒪pn�~|�Ԧ��t��:vD!��h� ܗz��G� =�=���Z��hZ���C�3��	�㊰�r�B��R6`.�C2YK����wH	%����Cg1�����$$YԔ,� 
�l�=�f�xB=ƒh%�4H���_����y�X�U��kO./�w�<�����w�Z}����K�����&���	⻒�&b����^����;2	�ދF�}
�v�E����y��f�-�!����d�vt��al�ݮ"=n��'��X-C�"RB���e�)�A�X�'�_�?)f5K� X؄�^�a���FͿckZ���+��X� H�p�a�u��`A�����MD1�Fƣ�M������ˠ��;p�s�&b�EK_��?����]z�u�ߋ=3���p9�Ξ�����g,D��q~�T�D.��Q�D��M��V�Nd��;-}�g��.t���J�����s��S���6�.)g�M��7��Z��#O��)�/Ȗ3�D��{�j�f�jw�)�Po�U��ET�ib������<��^��VB���wW�5��a�4�N��?�?��$�a␲���V��p3��[z��=o�Nu�Ѵӛz��TNO}Fc���i�`�v�v�����B����_KQ�����	�pb('���s���|m^-�-{��۽@eX�����x�Rf*b�j�cz�RY�9�9��8�>:��&0U�h��C*�Ze��?� KV���u���+�7�H#�z;�*NY��"��%>^l0-C�����k��]R&���(R]p�yZ
p����S^f�9\���H���E����ʻa����LǢ���"%mjℐ�����*s�O���7�i���+�A����~x���ܹ�Vx� �w�q��4<�]Ʉ^P�$f}���M�eSb���^Q�U��?��q��R��{5���,]3�]�����g+m�鶿��vV����(7���Jީ�S
s+_D�#�Rz�#��PG���e�^/u��x~ 읺}4��l��^���"����3��q��XR*��M�53�*Я�)G�,mU��(᲋������$���-�R�t����1U�AX��ą{bʂ�p��A&\���?�O�]��c_���JnN#S����� E ��I�{�)u70��F-��[��;j����~ŭb�#o��@���AZR��J����7c2=�>�����S�����DGl�X;0s����*�?1ߋe�����\��7�;�p �4�$�»J�?�u��d��9 ���wm�1�!C|Q
���6	��8�#�t�[
\0�>�������G� v��~��]:-o�{ItK�<��x�����hؽ
���dWK��?�G�H�R��Fa�� ,��ߓ=.w*(��M�h^��$����Z5	S�^i�Kg]�1l��@���g�������s�������C�\m�����;���7��j�N�Zv�5��Y�QV''*Z/Ipg���m�B.Z]�h�c��|f�(��t�DϚj���d�?v#%M��bj �7����!�v��&`��Iݓ�V�&����|y�r�0v����>�� 3J|��xK��^nn�$���s���t"@l��ǧ~�>6%O�/<���ջ����;�ߵk�w��W���b�Q���P����x���2E�C���v�=�-��zm����3�05���`����#/�
�������퀙<�5>�J�]���@�+=��G <�ba��喳�&���[�+c��];Ģc���	4�F(�^�Q�V��vҹJȉ_��Hh���כ�$����L�m�;3�ͭ5����t���U�S{ؗ���ԡ���ꗟ��>����*a��Ey���x��Ō`&8�7>!�=��GQģ�n��Q��:T�I`�ks�!����(����,��gQ�T���B�Y��^A�J/-��L�!�e�*\l���E�=M9���!�͉���	�$�v2�~�D�Ɏ���_&���3%�݁UW�+���&�*����� =7~�jXVS�U�� ȒYj�b�7-S%6��1��A��
�V�r����1��Bu$���?�@4�?���8��^Ϲ]�+��Wʶ��_9I�_�0Ѽ�:�� �4:�>�z�a#Bz�wo�����L��l��L��$�e\|kVg��Tm�֮��ܵ�m�6K��C�g����8�K���:Cz�ה�[�;���b=z <��%�W��b�����E\R2Em8X|�z��q���xs8�~c���M?۔x����-Ղ��0N3~�EOp�:�<]���T�p����%ӂɁ6���G6��F�?�j[�ȝ���k��3f����6�U����^:Pz�������^���c�z^7o���=o��|�G���`p�2�0���%)���[-�)��*p�� Q�g�H� ���W��qSl��,��\_C0V�uD���g�-��� �?yE�>M�H{緁����ʵ���_�e�m�!�8�7����Os$9&1�V��+U$ywQ(�/�tvc�,$�|r`�a��bc��	z9���K{D�C��=mj�i�X7����'[q뿰����iWo�V�ӝf_T]Hg`��d-waa�"��yۂV�cΩY-�f�2p<�����q1���;��+f�~�+r�Ng6��|g%�6�(��Vo#d�V���̊�vV�(�����?ޱ;���l��^�}�?%ē�	!�ɳ���E��ǒ��e���˟�u�M�9����=�ن�zB�񇓭y�j(&#Ѡ���3a��U�l}b���pYh�|���y��D\b�xiR2/ �άMy��J�l���� �����3 �{ɳ'��6N�@ƙ�O>H#	j�p<�C�`(���d��I�V�E�vR�Ga���rI��脿{gn�ܿbZ��d�/����)i"v%I��!"QZ��v Yob8\쫏]���b�	K&�^�RN/+�`��ks�d� F3Q%���ͬ��y4�58��-�+�C�'�\D�ۻ��eK��w�^ {��D��p5��W��
��L	�ہ�����M�s�%��KǰѩB�*��/{� �.d�.�F'U΅$ֽ|�g�g�C.���pʚ��g`���z߹�<_X�� ^���Ncq>�$W\���3�v�"+�"e���h!h�+t+%p4�ր��_�Õ��Ta��s�<\����]_t�ե�{�A����+�5/���L�����3�Lw�l���x�Vgc��S�Z�\�����O���"�J/����/�e�Z�\��sWHt�B�7TtOo�O���	�3vS)G���,*�Nesz����>�?\t~��RqQ"���f��L�8�� �E�i��7T�ޑ�/�^�:�0�t�o@�4(A�%��Q�'֌����'�o��Q�$ѩpd� �R�ГϞ�_�v�15���V-��ܣ(T�����!L�\�)l�$�3NǸUf\՜�u�<�:�4���3�Gc]>�qZ�D���4iE�,�<�줌?�FV�{��ٜ5hπ2}�׻��F��ѶN�%3��y
pMV��e��+�%C.��	��|���X?b�-B<ұ��u2y{pʔ���N�en;��P��X��`1����g��=��դ;%�\4�B$:CUP®���;�e�e�"�ݏΘw��࠮�Ұ�M��M�m�Q��	? ��o�O�\��ce�qҵ�ۺ��Z�a�Չ
���5l.;M�F��4�ӵP7�ti��}FÍ�����Z��5:��`�����B=�HO(Pi'��e�&|���ǭ[r��R43Ыcz��"������8d;M���0&���WIC(�<�t�yv���xw��+��v���Ĳ)��&h�Q�H�P��t���dA����`"&v��q�N^a�I�}60U�pۘ����w�g8�٦ˌ��}����*�[�X�vlÊAC�1B�͘1�]�x$��Ж���!RI
��W�,$��.�J쓭����FJzI!��M|�Ȟ�Nh�gf�=�Ǝ-l��g7���k�X/�0;�or_����x�6�NQa���S�!u�4�q�����1~��r?���H�]����kh��Q<�V�g����}"���ل��ˈ� � ��%ěG��q���;)S܀�P��M�����뫯%	J��1ڏ��GM�O��5�V��,0x���D�,o�5�*��X�����z������ֺ���:ou�1qFQO�EA�jv=��{b�f2P@,�C4��
���G�՟��}Kuйa���#���Y�&'>#=������[9)�~XOm�zZ~�C��ϊv��Cv�s��R�pH#�[	l�OZ[���3�`�]����Vy~�8���O��]KԜ��l��$������*(:]�-�|6ې�}�"�v�2��d�4�zYA��=�(�fdOU����&OG�E��>��Ꟗ�z�f��/R����_ġ�m����%71�p�a�ӯy�uιY�fţ���p��ky���*FL>�����|�F�S�>���?�r�ʨx�����} �
�y9C_	���b��	�p7 �HyLK�V���k���:Z���Կ(���]F���	�-����D�������R�G�%�i�7F��qz���ؐ�˟�/�������K� j��G�'�M&;C�,Wޗ�k�|6{g1��2�G��b� m�J���(欫�/�`\�$Ρ��t�z��Zj�7?y����їtr,3�}�9��R\�!���(�u�S� ���QkMS���r�>�<��8��C��J+��\�{����e����< 4:Ix�~Tw���^�Ҫ�Ӫ"���Z�E�YG@u�4�Lt����SN-a�6��G��(C���6t𲆵�K=8[�E�^$�v ��}�'���'ז	L�+!=��:����8/�z.�iBU��sY���d�Rk.��@��	we[�ه#T(���bФ��.�����`��l��4S�\�Nn� �W,�n�ɏEb6jּŬ>��e�|�V�L)�6MY*Mg�e��b_��L^�=����I���rᖐ�t������q��@5�^A����
↉�=�Y ּ�h��]/{Ec��/�]���=���/NvG.B��	����17ϼ�bm��ݗ�G��5�w%6ˋ̿K���~�cQ,Ȳ	�$�m�|�d,$�� C��fo�`�Ay�[S����A�4B.	��.���h�(�Zy6Լ#o�N��G+*�:hR�[N�"� -��:�����gt��橱���	��iQ�ѹe��N?��w�6�����c	�#�y�f����Q����� %`rłfP�F(t��*e����x��j��M����O/����	oO��Ta�~8س���W�0� ��Gv5���Fb:n�Z��g��b�)��$�� �H*"�TC�6��l6�:z𽆄Bb��` ��z�x�d��6�m���X�[�O��B���
��K���$�k�۶��p��2�p"�yj�;t����S�a(���[��@�w5_�(��
&f�o�a��yUn7?�$}��^���)oݚ�vFø6�j*��;��?i\,r���u�j�6����32>�;�}���*�����_�翬�.Dp�s|nIPUdwA�q�*A���}�!g�O�!�	���d�d�����m���u�:lSP���	�D�LBi�2�3Qw���am���P�7{(}W��kj�Za�y#�/�,�{i/Ղ�Yp�7O�@�*��C:o�6N�=�9|��S5���ʙ�N��ꓙ����0��/mg�$�K�������#W����k���1d^^�1g�M2X�Z��D���A�����3� ����H��ў���+���#�;��4y�v<8!��j�kG����"H���e9�L뽐�8Z�v=E�h�uWE��Gi�^�^5��P�`��pj������9���r4Y�Ή`A`��B�����Z�63COV���8܁�P�7��Q�����T�8�7�z5���Lr]��O|�h�|�D�FE7aH���| 	��J-�����r�>���H�K2<��>����������mk7u�C�z�/����a��|Y��j2�Z{J@��t�0��)���O+�.�1޲]��M���&O,�#^1���.�0�44)і��Id{�
ט*�R;[){�bS�_�-]�JT�C\�T��ԕ�B�`�C�1'� ��ާƿ�r���72�[\��?[
9��ٓE,�LVP����8H�I9<Ꝇ\n2U�����F��D��䅺���"8�-QVh��ދl��c�a't�k��z2hj��b_:�<�Ф#>j	�