��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L���VFjU\|=Eʅ[�4��o��?�l'����:W���8�����$���������G��3�G9���wM�}�d�� �0ۘW��g�F%��O`�l�u��(#E��s��[33�v, �ؔaf|����D��v�JK��y1����̣ʱ�Mޥ|^}y�`=U\[o�ۑd,`��pg3��Xe������>R�8��K���]����l�vLe��C.$s���V�D��3���K�h�5n�Ä��p)7Iy/�����C���-�^ɾ��Mw��?V��3����~yZ�i�c�9F�'��dX�����^Q��PtMɗ\$�T�26�D3S����qx�c��͂<ѝX�Z��F�DY�'���ަEM�"(�g����`��5�J%Uw��3v��N�*6������
&�CF:�2�O�蠗S۫d�?=��|��K�({���7G�G�*r����_�A�/~���l�7O��a�Kk��� ՞��@���t�,a��0/�0ޙi�1�i���匶�f�F�Y�E5��-�-'F�PԘg�@vʋ�"��V��e����+[��.�!N�'^���c�|8��P�`�xjh�������DL%�� �8�8n�f��l�c�����%:�ǑSd�Lh;��	��$�������%�E~�G�����b���"`���k��ͼA����0�n�@BI^`��gD	��|��::5�V��߇
E����,<�'?jk7�k	P�3L�=�2n�ʏ�n����ɷ��J(%�9x�E>6u��l��Ê�""�/�
�B��Z��2n;�ɇ*~3�u�q'Z�m�ѹ�΍,�7)��Hz�3~Ub����	�J�<J����m*F����*?��ɔ9�=���u]꾫))��_���x��91^�p| �h���.��
����j�K�����'�����V�G ��ٗ��vv�����4�Q���=�]�]�#���ɕ8��T���)��<�WT~D~S�9�)��_Y��'�k�xwE
�3:�$�t�WF��#+q>�����_vZ���Q�`���qf�PDרU�(6Oa������-Ɠ�|-�x��c{��Y���!��%�g�ki�}�{�����N}�\cm[^p�{�
x\ɘ�^��&�̊��H��4����Th�&?lh*	�6�: J1a�EJs�q2���������O!Cޜ�jԛ9M�5��WI�liU.5b�,����F�E��{R�"�1�a������^��ZH��RW��ruh��iDhÿ��Y�E��_+���&��I .�P<���:�Př5Tǟe�b�l���QF>�ίf�Y���!�~�����9?&R�����ʟ�J6�H���,���l��۔S�D囍@�P�{����<X�/�@
)>az�(E�Ҕư\�o�
��ǈxF\�ު�4����Ϊ���E��/�r��q~��A����k���nh9ɥ�2\aØ�9ԟId�P����8�#��J���ڨFu:�~5N����|@�D5K������9ߟ>�L'%�S�{�(ƪ�6q�j
ٝ�Jm*�M�֔�4:���T�Y��͉�/�[!VN����I8���y����.�k�EG`ǒ]�I�Xۏm�0�{�`[*�D����^묦�P�����l6�o[�\�8r⹬����[�f���c�n�g,XP�T��޷�"�\=��nV/GqJ� �$�~�v	��o�C��PiS��c	����;;��L�hni+�&A���D_#6C|3��{�j7w���P��#.3����ў(�CMi��P���hk;cD"_�\��B��E�6���]\�����^���� �.����g:��gA0����pm��3H�Dk[ÇB��Ӗ7�	=�O�5�<���?��=w�s�C���'��ҵT��x���%*�z?��ϖ�i�7iB�ص�|֡�J�p�}^�K�t]�l�/5���9����1iM?EU�Q���s�/��]!F���.v�� RQ�,����Mp"��'����$)Yuw��E���խ����\@aK��*�<�Z��N�9ӟ��W�����U	�k��mJ;ޮ���jN���YO`��!:'�k�ȟ��8�1Z���$+2bB �>9V&^a��~0E�4<n�g=6!!��^���ǣ���:�53�g�S*��F)�[Jy�N`òQ_�uA�kg�zƘj�nw9�+~>0V�/�{���S���'S2�ܻ�g��_p0�f�9�({��S};ۏ\�ѵ	��I��?	���*q���_(L����D���	Avir�~]�l��`<D����i6��k֪E��)|
��笆s`^������$(}���y �@��Em���m�����	u��=�Jŗ	6Bb��
&k S���H�,>�j�ng�8K~�;.xdo�-��תX���s���L��=�/M�O���R5�)k�����O� ;������yk���;��WT����}����sC�g|(QJ��?/�������8s&i��E�a��K�C�l��D�cs�d�4LV;M}� ��Z*6�^��/iF��i�$��D����b�L�{h�!$B�
�+6;��\�B����G��u�ԍ�ӫ��?I��ӭ3�C�^�9� �l�w�/�3�Ʀ�;�m�
�~Z[����Y4����T��=�ۍ���J6P��>��
�#[�,�ac;�8��k�w�9.T������M�Fn�сf$���B����ż ��+�[��l�r�]�ISE����6���	�˞�y���w�5�9�y:�h��q}zb��p�^�&�2SGe��Å�X��eA��N���GVi|6;_��F�QS��
�W������	4�s'��ם��"�.��/��@b)%�-f|u�b��H�^�n�QU P���D���8ֵ�N4�M�=�{�v�����/�D��%���;$1��s��i"6Z��-� ��l�=��p��ʈ��!�8	vlKR/�	<t�HC,�)�|����T���Ԏ�Q8`.�a�ڍ�[o08*����P��e�>^�!3(
[�)O��YX��W�UӐ��d�Tw"�|;am�r#������5{��1�۪�}�CX�b���>T����r�^*��/��p�h޸�R��WLG4ѧ�Y�m�|�<"ģ�N��m��M18���Y�˂�L��dJ����A4���@Lf&2l[������N��S?S*��?@�~;$�1Zm���;N�����նf$)�Q���,��\��n��K;�B>��u���!u��F�k�i�؜�o�?A�#���V�ާ�u�08�������#��ƭ�EA�Z�=?sxU�����[Z;<���	�������D���=��	@(��9�uTYO�L������mw�s�f(��7�|�m��a솉?s����;����1��ey��Nq�v�?a27�9>&�b�E>�pb�PԢx+f<����!�>(6pb�p�C�����ɬM��	/C&�:X�E�re\+	�P��?*F�O���1��Y퍗vÐ7Q'3��}�%�*`*�,2��px�[��ˁ�H���̹Q�aڹ0��w��ɚ�u,�I�]�V�Y�d��-�fL�]E,�����Da���`�����;������ε$�âB�pҖ'2 o1���`S���e�~��&�#`�@n|��s�*`��ՙ�@�Z���J&�QCN���wk��W�3�Oi�)�t2�QO���
�E7�r�v�FՋ�����	�Ԋ����J�
�Na��۠�*ۀ��(F@IY��^�6��\v�dZ���h�F��5�u�\͓f�H��󈗈�ש�J�c�@_�gk�~��, �����}��~��� 2�!xS��R��'qlZ�V��\,��{�
QP<��o�sVg��Zk�{c��:��ECuǾ��u�U�@x��e,<	��^�Z�ʀ����׍�U�>
l�A;{}�y������
;SPUQ`(�jW�j��piZ��U|J�� �����R8[q|���wtw���.��#"J�м�u��/f��9WT�07�F�E�{�Q�M�4�߻���䩁x��)$&-�����$�9n���{js>bۺ8�_^���V��`#���I:�j��3*U����O��a-"�VYfz�E�!��Y�V�9�5�t�t�cS:���B�}�Q������<7��"ht��
4'�q��ݠ�?&���̨b@T�J�����v^�|d�򝌗�;��қ�����3BS�k�W�22bJ~��m��ݡl�CkA�����4z��1��N���8���x��m�K�|�~��Yti�C_�סsY�1 3�e�l�
;���wA�_Q���SD�J!��;ұ�]�|��8qa_W�("��VͶF���5��|7ne�jq�gm�`�ZE]��6fJ��RnÑ#���={c�_{�Nj7�| m�;�
yW�9tɾJ}��v�$j���5�v���r*q��xy-x�Yk�e�]^�$���)��".�!����@�e�d�]80',c\�zK+�S�F�Y��;/Su0Zo��zJ:o=���P�!�k}*:RL�������.aS�K�[~�V�w�d�������"[Y΢˗ЇD0 �^��W��f���2��{l�px�8�N�O��˸l�#�y kw�cW쀺�M�i_@nn�߀!.AY934wTQ�����R
��PP,xa�ʑ�<&�D�����C�ނw�:�s���mA'U2���Z�E\o�	 ��a��K�Z]$��{���R3���ah��i��	��l�GF��S��U�a�k����X�U�B=�P���8:S`wѿ#t������޵�vuXl�yB�_	kX�?��D�|�?���/�ɾ��R����MZ��z<�A�8�Mb.<A�qBNG ��㇚Hn:L��s?���I�㢝�Sd��CNi
<���2��<hD����EK4Ѧ�*���y�^��N���#���ә���V��a ����5�����l~f�VTG�0��O�a3:������4�n���^e{>��!3K$�~U%2�9}���V���v+��ɇ��X_ꖃ�6h�^��.�z���R�	d
�{��	�W�}0Grq�_�  �+F
��2�(��1 w������or���b+� �o3Fkf-)�$v�&3�� �<����k �E�����J���r�Ć�6�EXL.R�z�c��)�jYY�)=����2`�$f��r������)�����կ���A��z +W�\�:�G�/^�$)!�U���]��^? ��@�-��a��6�b��<rt�a׶f�����)�?�!7]3Ě@v6\r��5{���1����W�k���T��-_n�a��s��ф���i6�Z!TS�9Ԋ8yw�; �%a|s�L�U�j=��R$�6}��,��n�.$��� w�d�%t$:����w�:GtS����	�(s�MR#o�T$��٧A��M��/z��Fs,��}�n�P%8vbm��.Kz��]J��}�e�Icq*�o)x.hU,�F37��L:'�&Q�9�
��T�bT&S�ȁE�C���=*҂,W�[�d5}��5��'@|58d��N�n��AHxHa��	���A��:���ly����[�-�fA�P�w�������
�|K벚�&��<\�?	�M�U��<<7d_����.�I��眍��_�a�r���4��ǻx��!Ơ��-��r�x�+�e&%�H���I�m�CE�{�� �cY/����`#�p����-aq+�1������{��D����4����)�s�lk
�����h����G%�G�k}��8�ʞ��ݽk��_
��S�'���w�\#bn΋a~E�bln ����.Q�{�3�����,?ٸ)�ԓ�^k\v�X�a,/����`;k��,��s+�W&�9��n(�q$Ѷ����������o �e�����u�nQ�*~�?�A^`�q��0}�:d�u%D��q�]�n)EǛ�=n}��s{ t���q��z��d�MuK9(EPz������Z�u#.,^�e��Ї�����?���¤g;9���i	�ٙџfPX�BeU�\h�o9l��#�o�s3\�(]��ӌ44H���4�
W�%7=m빝M� �|ִ� k��wV���|��V�f��ӻ���	O��O���jeo�z����;{MsF^���)�&��C{:v�{���(J>f�A���8�h|�ݥ�8�]MR,���>���s+	�M���$�^�am��v!]�d��5�x�/v1�g
�2��Z��TvT�?�mo��Є�ep���q�ޮ����`]���B_��@�	���̫�Ė���_�I<#���Dxhg͘����B��a:W��'�?�O|���ZP׵"�o؅�hN���';����B��Mp"~��"!�Yt0���<�G�9�AQbH"���z�^���?�N��!�nZ���p��7���Yr�'��H\شe��>:9f�aL�˞��g>�Mo9;;�����Ai8t{��;\��V�b����]�8��3\v&> ��N����$ N��DuOKP�V�	L:��`<�>�^��q/w5P���-nq�*"wN��ﯵn����f񩽚��6����џ"L-�B#������Wy^Й6�oO�:PKZ�8���|��u�^�0�@�Ɇ�6�Tr���(c3����V��re������	w��ۘ�ޮ1���s���*��x�.OE!�nh���oJ�K�L��~�������:��g8r��E�f�@ae�_U�ⴭ|���b߫᠝��u6��-�|x�|�-�n44R��2�1,_�-����z��
CǭW�)ޘ�>v#Z^AA6!X���V;���\�!�`:S�Z"�r�cv�~�������v{�0�ݮ?�q��"��L�M�*�Һw�;^��l���.�I�r�s:�hOQ{�S�ħ��ߪ����l��	�<p��gN��be��T|��Ậʘ�}�lѧ0q�&x*��bH��'mP!��� ��X;ס2�G���T���"�Ԑ?��R�6��O���#�a�:F��X��rj1���?^yu�b�_R]q��<K�� v2���I�H"��;|%�S_L��Jt��6��^�vH�ߺI���� \.�F�x�uͰn�$ݽ����DI���=�b�n��bE��k�\"�&�\k�)sz]5���.�1J���� ,�x��L<�I>8�V������E��d�Gk5��Sd��3���/�L̆>hiS��`�:�ơ����񵨜�������%��@XZ�-��7%�)�܎�����c� (\�+-�ow�PCX3(7l\O��'h�U�y@ے�^����/�'����A��f� �^%^�dF�"⮰���0�����;���}<��(�T%[�o�@�����W���o�z�*,;�#���P7���did����; ���k��o��{Of6�vj7VQX9-XQ5A�c�^�N�����!(�0�ǭ��f�� <�&�v���_��Ģ�aYp��W&��N���[�ĩC?@Ų���Y�p�2��5@?($�ٲ <��x��1���fO��Io�eb��Cw�m#�Z� ����#��P�����^��
^:�Zi�Gb׎��if���@�����6==�	�Tl��O5���E+�#��{�$kL1 x��h^���\����k��C�F=�u +i�1�����}�˛AH�ז��U���s��R����^hB�^/�xe�&VK����쵐j�C�L�)��q�Q�|�5����t ��d�����.Pl!�������	�I7|ޠ���z��2�x��8 0me͸W�FB�Q[VW��4( :���S��l쫅`�V<�MA�]���_�NMe0�-����CG�Cɳ���d,8�ҫ��5.-���s�*T:��5�F��n��=@��y뵔N*��%�djD����$�ga��9���Z+y(~փ��n z�i��i�S�����c{��s��K�yM��(��	���q�f7|)j(ri�Cn8�3qS�����
��-'�v�3���,�%SO:P�]��&Mb1YO �F�wF�;��nBLl�H��0��
��No�:犯�+# �{��4=����X������CTTF}82�W1����+M�����W]�����qI��h�@�&�`9�pB��%%����S5��
] q:������四�{<��<�>`�鱛C��>�Gs�n�d|&����.�'��L4��2U��@2?F�2���h�#��+ͫ��*}^+.{CaX���syIr�]�xL�O�(�2N����˽ F�Rh�m�����;�l���t��P��K���C��NIn�Ms]�˱&�#�9K�sI(��-W�d4C��vňw&���g�GH��_qdң���T!]:�CQ��f�3�o�����i���ul����x�r���<�6��z�C��P���e�!9e�[@`�'�0������71���%�
��2�rxP�hF�y'�"�e�7�<���%�C�*��_;oT{�T���)1����+��W�y_.�k��؟�ނ�B�������z��X��n��E����\�"בT�	>!�b����΀JS����
���ڨ8���.������Y�#�������&/�g<�sa�)�y��:��\%���r��T�)���1�d�A%9��S!}j�4�|�6��6�gS�ă<��&�k=�i�Dܢ"DY����*ӚK��{GH�ߝR�5+wam��Abڊ:ƈF2�~@[H0����F���ra9������X��T	+�g)r0{�:���l/j����1����"����n�I��U��/Od�+k.�X��h��f���:�Z�"(�7���]�F��������(���z/��2z�<������E����TͿ&���ㅱ�pNFe�&���J��ՏsD?`��C�gA���$�6���D��)a��`ߘ��3�, �gp֛,�b���F	��`]m2�g�|+����أ؎��S�v�����
5n�c�꥾�eg�Ҥ�S֬��u��$39�&R(j��l���a]z֧h��tȼ��z�zlTVBs�	�IͶw�t��7?�3a����v���s�D��Ią� �v��+����c�
D�޷��g�w��D�pR��M98��F���~���Dѿ�3�\mC�	2����&G�a�+I
9œ�� ���ŤQC��ޟ�>3A��N.q�1�����}!�+�0[�dz����8��A�1ڎ@h�:V�J�nq�$����k\��*=2�볡�=yǴ�*��0����u�ۻʹ���]m>M���`N���7Cp�g	�g���Y��.����+Q�Vo/"l&0�/?u5w>�/)R��岱ŬM�5�Љ&F�.�,�텶SLڢE�o�*.ۦ��]�!T/�wn�rmB�#�Ղki�U�l� ������07rZ�����I����2,�|Oܔ���LԒ	!0���N77�͔%��@\�A�,5)2fd�-�GH[��#)6�&�Ԗ>ii�ʘ[$�%㤎�R-C,Zo>2�V���2�B��.0�"}�k�E��oU�f.4͙���^
b���0)I;�=��/R�_��G˔��Ι�Ŕ���d�E�~~E�槠�H+�D\O1�2���B�"ʾ�
�kQ�vgd<B)�G��R�ٗg����3ƌi�L�l�(e�o��G*����iWL>�`����y����4�vߙX���R�v�f��5��	mWۣF�1��U���9�w����I�����=�@iV�2���>P�T��11�^�4ֈ��䒉k7}�<�W�ւ���ą��1)/�����~}���k��O���͠�?��܀�,�]���㖕�2m)9q��H����H��2�@�!H�˔�i�����e�e��=���ES����Ȉǰ��=O/��$�O5��d|��iXU�A�[���L�<.i�?����β�J����Sc>g^8z�_�m��2��q��A��5�q�G���7�����;u �6����:��}�s	w舎ZK.3R,��C���t今�0��������1� ����a`>cz��#V�d�ci�/`����݈a�G��mA�F���f��X	���r�*P7����`��t��� ��٪@� ��˫O�R����w���nQٮ��#��_(�Z-<u��.�����.�Q�3�sf�J�9C&L����?}�.�\�C��aA,��1�	|�e��?�s� �+s�!Ս������/ذ��&������Gص􇯔��;� ��u/$T3�j���TgC�Ʈa %�ҋ5ŕD�R~J�q� ڂ���n�{��6t�w������w�cHb�=��H{#�W]�C�N�8P ��+��ge\O�۳�nq�z}����U&h�*�`�C�6���v�o?��9�r��j�	�a�"���]�[1Q����/���z����iS���o��(�3ڜ|�����p�
��o��oVK��s��6;�f|dV"a@��*+2��+�`j�[�Ra<���?X�b?I~�;7c��N8��0<q����_6f���\8�m�����Wx!�G8���˴�3��C����m�s{��h}��5~����p�½��|�|��[1���([����p���CФ�vY��V��7FbA���*�͘�͋�WQuq2h�L���O��]��RTh"�������A�	F���=��"j��g��R�r��*mvY?��le�>!``1�`&�s��F����ro	&M�{��a�6�7��|4��/�8Dj��O�xV�"��yq�PcN�گ-
��}�Π:�j�f�4E �A� @x��~���c)��G�����F�/XBs}˵��c�[�A��7>2�پ�!lMjmaiݬ�-RK�1��޴����������Ϸ��R��#ōg��S�f��nƜk���ܪc>ה��
8$|�����G�Bx���������Pu�ip��Y�?�hI]��Y�&�^�t���a�j�{���R�{&e8��Ｗ�g��h�`c^�Ck�ʨa@t`�ngXB
�_ο+�k�/_��6yp�;�����=dS0&���ߤ����j<�83��1����j���d�Lʟގ߃�K=%`2�:�4��@-���=h�ec���Ak�j��\�Q���z�� 6�-��0��_ ��;�<��ņ�>�voX�Q2�)�ݡT�/���/�!S+��k�A��?J�v&�%�!vZ��r��_w�C�(��bd�p���{�{�KX1$�_ҿ��%��W���7��5����gA��E�@#��E�M�� (o�Ը��M����AV�2�Y5����[�=�_�q����wpt-eƴ��LO�W���🕕{��n��ȢO��pT�/`�Z����~��f���^-�F���Iz� [iȡb��CP�]1i�3���=/�ϛt����S-޸��������M��Q���r�[�g�7�����&1��S�1�$��(�pI��? &�z�/*����(����������M�X�@��������Z�D�g�O߆.���U[<9T�Y`N�e&���Y>ʞS�GQ�`��1z�cD��X��DԖ~���DIbEs�%s~D\1����u;��ω03.v��w�4�� �+�D�P�Z��*Zx���r��~��m�q[Tn�ՐB���e�I���<d"B�+1�*MF�>R���[U���gly�"��'a��,�F$0��L(1O��;��o3]AN���Wb)��\�O��٤s��j��Wl���ɶE���;p��0LW�6�$��3���I�/Mi�N+���<����ޯ����S���6{ҕH���I ���)��p }�u5H�|�]?��_����&a�iz���9��(���$7�@�M���@����^�����]/2���.b���k������������$���βI^'�1�/6�ܰ͟b������p.��|b%fs�WX��br�hhASy�q�&f$̀P���-�̟S_4��F����R��"�>#V�J�S9ك�R{�yVS�-�[�! T\+�8�
��l�Y�T��Y�����J���!��U=�tg� �㯞kG��2��ݝ��r�c8�,>���ѝ�t_z�-=��-=l�Z���S6T������ʞr8ߠC !N��	J֝q:l�<̀�f��	U������C�#�i�B�sMc���c �Fn����2��5�Y'ߴ?�_�S���Ϻ�ـ�'$m#O��j��7O2�r��Nخ��#�����H^�w���}%q'��c|C�{�p%�d���65&+`�#�"�K�������4
~_��i�x��XKIϯT-�0>&4S</Y:���ȓAZn��T��w~�NN.��:���N?�U��A��6�(�J�B��Ϧ�K$E������is�THX}�������A0��	?	L�/��Eyӄ���5�3��i��;Ivr�AP��b�_��7.'.+PM�������ݒɾ�^�BKƜ5�<��@����o3V�
,r��b{ɮ���h-�_-��`��TT�?��ǈ��H���9��1� ��&�jVt�$U�xm�h�N�A��Ɓh+��e��@k���T>L}�Zm���:���Vw�RtYD���DnQ���	�R�K�.��,>��W[ڬ�`��K��!Do_��r���Ao܅�w���|�Kp�`��tE{�y~��"��ޑ7��m�)�P�,��S��Mk���4x�/d���9�=�՜�k��Ӹ���=�Q��eeD��]]>�q��6 򘲋�k�t�$`#Di���i$��T������թ ]�G�jA�p�T�S������|"�F�d�������F�H��L���m�z�`%���7�
r L���]�_�7ĜՆ���ї�eྻ�=\>�M�͸r��%�\�+b�h-ᔌ�΀[��Y[���'�.�[�W7R�ܢ��ݲ]�t�=�B���������Y�i�d���L^m��أ4\b�6>s�e"_,�F*s�{��Ɛ*
W^�����
�>���E���@X���a�8+u ����(9����R6mV~����:Zޑ�E2�Rs��6����Aa�W�+��TI9��
ߢ�PmD�:�cx��]8�.6Hb%:�S��F]�ZTn�_�F���k�Q����P]����=�t�mn�A^36�8**M���
j\��9g̑�d��˱��$�[�)�3��ͩ]Z�ִ��џ>�`c'��D��'�t	R.�6�ӎ��D-g�8�M�!Vz�� Ɔ
�(a��8S"~�9��� �1U�te��g�c7ƊE�g��.��S��+6�A�9�Z���5^���>�U~�Ȳ�=K����d�aw�lX$����}�BYW�>Z-�ȱɁ�ْəaܡ��K�ß�����jk[�<��������__�xk�*VHb���{��v�*�H2�ڝ�	G��8ԈR�P[?Wt�i�BB��q~9�^�d�)���kǳ@�5�o��F)M�&+<�F�O�ݻl1�i3nZ�k�]׿5��=������(~:�/�ۥ<W}\���Y_Ou�s'y|�l��a�)Ƅ28��+&��Q�2<�� #�RGmd�[_7�M���԰�A��Z|���p��D�PxǨ�D*լ�cM�����g�el"�f/vi��'��ؒ�l+����]�����P����Ln����d��i>C��Tm՛�#��+��TF������'��P��n����{(g'f�_z���Lp��Ř�Q�5�-~���b�x����=�ޔ�9)B���meI��|��Ɗ`h̼��
���^�6()a���p�ٙ��
�)h9����*EOB@�^���Z�d�b������m�;"r5�e��f��Ěi�He�)w�5�n�)���!�H0r���;�D(�����I��@̕�Y��R*:���� ������1
��M��:��
 $d"J�^\q�($_ǲ:h��t�ѯ|�N��|�L�Si�N���*�?��]`C����1�do�������'A����MTcUF����&&��80���;���ђ~�Ps� �zf�@�u������i�q�t_�7���®[9�բ�q?�} W{� ���<n����Uc�ԹE?�����9�-�EjҾs��ԥu�Z9T}�Rqs9م��`�]#�0���@�HLj���^�$G��؍�K5�8d��8�,�<��\����wp���e�c�O�ʧh"%�ߔ����Q�h{3��9�${�h�g�����>9�R�������w
�/�w�c���X�#*���G���	h~���$�>��I[Ƅ;��
F�[�n*�u��`
�;�3�B��V�H�{�\����R$��*Ҝ׶�޵�>�QO�o>��+5r@FK�	�}�8V Ԧeo��Ps�I d�%Q���.яz�0r2��xH	H�UD��m6'nT�nF�6�vy��=ؔ���
GW>�Qz~-xL���G�eH7�:	L���������T�tD#�I�M�0��e=F��P���!S����]�tf�e�Zt��V�!��(�$�2�Bd���b���j��(�w��y�74���������;��r�'Y�wrn� ���2���ˉ�H��Q�:�<7��b�]�O����(����o( ^83qQ���(=�������rE�&q����K"
yQ�(3ʈXغ����t���W30��$Z��
�*�(͉�`��25T�T�Ɠ[��s��v�NO�y�Jd�n���.t���&��r:q"&��8~��ZȀ� w��im��,�)}��h}b�l�oosir�JU�M�J�.쟳�� ���.��b��pE��?�V.:���λ�_�vL1���[2E���1��2���}���i��`�E-��&�T���2x�.9�[��E�D��낝4�#pb��;&�='gJ v�b�T�) �x�l"����;н�$�y�R7�.2�ae� �h+�p�I�M��ל��2��m]�p�W���
{�J��W<�X�����k������.�o^Һ~X�|&��Z�Auș�@�?�Z3��W��(����B�0�}�KI��ݕ��'��룁�S��z"{$���У-;̎��+��j� v@֜�>�.3��*+��4��D'rH��h�R���]�%���^~�bեy��FA��[~^&���;��Q�T:�w1&�{�6�����"K�ؙ�����gs[�6����EL ��dʇ[�_��߹�7A��k�$6��mkqP�S��-x�V7����d�X�k}nE�U�v�����wS��!�4��CN���yL�G!n��&�%ĸEI�y�tB�aЛ�{_B�7L�h�]YՈ�Dl�{4�g���$"�����cƝ������m���J�@rr�rƻ�`Ohu �������I��[���gQ�QX(OYwN�o�`%���}G���+�+D�J1N���>�â�=�%]�t!�a�89��4�9��[:��.C��eD�h���wR�#�ղ.3��g� ۽�)m]P/��kb���+P=n�������H��K߮�Qo�X8bj*0������6����HIM�Xy�qP� Z`����򞣞�,�k��.�nC�]��?Vܢ�f��`�QH����t�$�6��0������;�(�Z=a����0c����h�r)�S}������5�!�8c�i)������MC�l<�	��ų_>q�L���������0bb�ՙ~�4�[F.C�I��x|��L�l9՘*����K�1T9�����b��G�OIZ��DNX�4&��x
a��O��|?"g���i�����gA�{hr�3��Fy�����{0MR�\-�X�[�Щ�V��}�=$����@��#}�0�r׊������m�~Y%�U=:t0�_MV��Mf-�U�����m�I��0z�
�0~��z�:��Eg��.&��<f�La�ċ���_���3TB�?�qaq�#e�m3��k$��J�Ƚl���p����>L�́� �-����J1��%�6����0�W�Pg�x�G'r������캈
�#5�B�l�i�8�ai7=q|p�~�%��z�3[��P]|BJ����6��k�@SM=˝�������J��U*5t!���TAi��ω��̿���/�t��D��mg\ɭ:��
��|Ft/�����3Xx޹U�i��v�k�:4�:%1�=��`�gB�c�:���UG���)���^R�k����oY��G���R9��z� Fg��(�����g�gƻ�؍���y�M����!�e�@ß���@� ������p;(�{��d�=Kթ�c�Emn7��&/w[�D��*�F[:5�!K��Y�xH�uM��Et�c	p��S�D*�t�{�#?�* _H��Ys��ғX��&ORe�!%��\'" �A���$GQ�e%���h���X����z�&3���g��R�:i���r�y����E�(kQ[RV��D=���ĕ��#�YZ���Д�I4�8|n�n��%F����*�ڄ��4[�2,:s_N�W���X�b'�8�5)Y�<��<�QC��{���kS����,4���l7�;���Gs�>?���qW̔-eG�4�\�W����P� ��y���O��hk�}n<�J���Zړ>�RuMO��f�N}\�͓�\�d N.��|ڍ����j�d����8�)��!��L��/U�+����RDp�S�b��턬*R���||fW�T��U��Mi#�]�!]��uZ��sFָ�&*X�U}�eJ�	\�&p��ԧ`ҷ� �	�������Wג�ET1�#��5�׳���	sR�y,� ��o�T�S�x"���@Z��K5����|G����t����2���`�	��xExZ4g�n@^�_� �Ym���ɀ�"�_Aw��%;%��WW0 �T��8mD�؄�:R�_0�Z�� Z���A��q��;�)��N����*���b�� 3�鈕i(���*;��Ȱ62Ú$_����Z�G����Ө{^�-Q�=��S�)Ԥ��LN�Y/\_#����]aǮ�~��1�G2����?�q�\~�n��V�X-�(=5.AzMk���m�eif3>���W�k�:*�p|mfs Ѳ��X��D4������jxں�^R��#h�s
�}u�W֪����V�X�ʣ����~���f�A���!�m��%u�Q�ک����	�
����{�۶Տ�b��7,	A��u����H���T����'0We��?����з��.�e���Xt�w�*�"�D��@t��ۚAz"��"��wӫ"j��	s�jvX,�'���{��֜ߪ)������{�N���VO�أ��{d��6���N�:"Y �"���� _`�<*�;h��K�r{M��Րat�Z�31�c��a�:	�Ԛ�������̩C�R�yh�z�K��2���4D}-#��Z@Ye�Ge��3B<�_�����Qcu �@�	-c�Ï'Za�	��pE�gp�@1�[�L=��Hv�,��;U����ܚ�\��:߬@B)���8��b�Az	�.�I����g�W�n�NK+��o���B�*~��v-E�C�s.X��ϡ�Z`�wt�n��V.� b����!��̻��WdKf�<v�9���2�]���Q~��7xB��WÜ�|����7h�%�~s�f����owA��5�X��¶�b�P0Fة<�~�l�=��1 �=�7����v��,) "����?�>�C!��	Z�u�>�Kt�VA}���U��5�ɟ�F�5|ğYK��L�T�=a��Dy��#&�m����9����z�����T:��*s�ȆR!0�"������Y�J�z���hK;��������fLe��ā3
��F^O']�o����?fED}��H�����V2��np٫p�*��LS;z��⻏�x<�^N
# �ǀ�����q�WTD��O �v"�AV���Z3�%����a�L3zP1��"���W� *͓~\E�^�S�n@:�����G�5�ޜ��rSW���^��S Nw'���>���Hۄ����N��K��G��S�3_��:��lz�9����d�>����o1�ٶ�	��-��Iɲל���^�@q�@:�Q���a�n���HqT��˼uֿ��!Z�t�;
���:�Sw�����,��}"qsp��+זU-�w�綪k���&�4�~���as`ɕ���r�&�wl���:*��bN������[y��%=��d�O�%�(I9`Y�Ra�m�ᑒ����	����#�4�����P(r����	��!���������?0D6�|�N�?�$,��m09P$�~k�{�Y�a�z\�<���?����r]���p4�X'�P�<U�xU��v2�c�PM��ʎ�%�a��B0˘[��mS}mg���F��P��d~�N�����u��]� ������b�B�$�l�Fe2�����Ƚ��<��*�V�>ڱ@��ؽ䊧�H�l4H)nAYLn�mļ��af�o&��#%	��ꛛ�q�2L�k���'4�,C�	�NӢ����M��Bѡ�_��}�A´�m*z�#�W����4�f3٢��T�A��`��5�򫬍E��߸(:U�'6�<2G��gU�{�BJ�$?��HB��ġ��n|�����7���TQOp�]�8�/�����8����Vc7,}��v� '-Bw�"אnE��wԟl�*�v)C�%.`Iz����7eQg�TջE�!:٘h$�]5uٽʌ��y����ϱ�bb��:oM\	Z��`���Iz'R-,����a�n����}4��Q]A�"bG]ܪ�Ct�ŵj�fF;�S�<y.	^A^�Y��^��?P�$�s���R�����5�^/c�2e9{�R�̌fn�O>K�ev��νШ� r�=�%�V`����w�_��3��5R�%͐��4C?�HHh�tL���g|�G�{�2:`(v��+�v���óп��qH�_�u����f�2�Ƥ'��$���d�X�;�PRD�����S�'hAX�湾oh�:o���S��L�^7��b�o��(y_�����T�2I.q~��i	��iN��X��^ߎ5��E�L4��f4T������j������95�"�ӂ�D��f�4۴eMhpIwF���?(���d��Xg}I����a!`N�Yz�b�I�S7>+�Xg	��I��p�g�0%�.2�b&e�����{������Q��XlԠ*��[��y;Pֱ$��{��Q/��5,b2�C�:rD�����pʸq'�3�}N�Ik�	hQ[N��Ow+�V`�U��od��>)��jb�k�1��`�&���)׳�nOʍ]�sSo�᱓7�����"ڇ3���h��k�z�γ�`�9��ˁ��Ա��a�V�)�ٿi��9%�srec�m z�X����Bѻ�2� ���U� ����?_��b<F���7�jc_��g+���#'����c?4��u�T��c�ڇ�:,�z��u�eM�Y�:ю��k)�RM,��;�T�|������a�~L��RT�,ޏf����-GBf��a�5��r$_Q��$A�1��t�f��(]��E\��cH�D�5�xl2쵄�d���*քN ���B/���C���}�bc���=�D22�W��	����?����ߒ-�4�JR����]-O\����@X��`}�J�ߩ��$s���%�C͓�}��g���̲�k�nm#R�#�2��)�K�����WT3n?��{���c׉]�I��]������ܕv�H�2�6�ZPa�<+CT��=���y�RA���v�[��8d"����}Zm�@h�������n긖(z�^���^�u�@?��=�d���/`�A�	XyDt(5]^A����W�'�s�i�τ������c����DK�B���/Ti!��dK��$��7�YF���c��@�IӂJC�C���~,�3d���w?~���KSP}ؙ�d�+���jȚ"�����Hԑ��%du�a�=���~�����@�Y��.�Ȏ׎u������x�����U��4w��&�_,���%ڞ�@�։\)Y$`T�0���:Q����:�9	Z��%�@�*^M��[��3Qd��"�E�Ol+�Z�n�, ���d�ڍw�IU�Z�;G�ђcN}����ȇ�tM��O�����܉.YU��R��]��ÞM#U�>Kqޯ 햯���i��\A������vEiN.��E�{��2]���-H�Bf�H@�ڐՃL��批�v9��������{<�Y�&���'Z%�7J�We��q�O���x2�$"�C��.�����'�>
K,9���kN�i�/=)��֙��ճ�r"tQ�%TN$��)]�F�|��R��fR>�|�ꫡ�Q��� �����lm���J�Uv���s	��4��>M����ZA�+c1�*z?���xɄ�#ϑk��=xaU����C���al���$�d[g�B�Q�\�a�
��0d'��e���s�=��QC�DWXش����O-y��{7����`rQx���7���I`z�*��'�#�ə(���)�	s���Y��"G�eU��|(:s�����yp�l��UYyE.�۱6�Č�v�V��Y=:T���'⹿��9��Z$�t��b��q@:ddw��zC��8����7f��Ҳ�!VV��	#�}` �1�P����	?�i1R�2�@��nؕ�ɦ�c�B����7$zqE <�OZ�>�q�꧋B;艿ÿ٬Onui��<���=�����R8F{:^����ry�(�+��o�~�ѳ��!������T��/'�y4S����ς�ʆѻ{�}�f�lQX]^0L�d�Zy�?�����>�j]�gz�5*~�ny[���V��R�I=�-w'�5N��9��r=�4��\�Rg9>@�	��vR��9���+Sr�iNaJ��a�7Q��yLǆ����|���&�MਙW����ՠ�����r��:���+�BF3���l�=/>]�?{ؖ�U:�LW*�<-�C
.�rs4[3UѦC��2\�jh��.�s���0��w�%����Z�i6�3��3�B4evBf�F<K[1�k\��Z��~$���i�+��Ч
�F�4���]�WХT��g���ێw�Dk2�
�鉡wIˣ�'��S�$.�)�-7���F�����3�O�\&[����v�D�԰���I�^������8��@L���5����f8�v��ܞS��!o?���h�3�\JL����G�~�
��/�r4��r�fe�J��?f��&>����v�8��J�D��������S2YO1ݖUqkM[��Ɔ�EfumXIKT;�O�$�:jë]��͋�Aµ1[����(P!���T�!�P+μdu�<j�5���>-�	��
�]����ަ�������"�YA���g>�%�T����D /b�]�񐐐�,��`�Jm��n�N�����d65A����zj���gK?�a����6�c��bk������#��:��h"V%������V(���7(&l&�`]��#��ʦ>���|������Y������� "�F�<��<�����p���
��R��+	s������Q4�.W�x�SCQ�ǵp|�������KfvKe<I����H����S�Z���w8���?"&���#��_��܄<���4g�_h5��GӦ7`� ��7ڿ�1NI��M݀7��}*j��Ԍl���؆��0�r�`�[DWU�z�Le!_�KȰ�t�b?~�1u񔦌a���vm0�K��t�vƤ�������gS(I�7iv��N�h0wd�w�m�Ԉ>ekO��R�.�`"P�E������s�
����O�H,R{���P/�=BW��sl��w���?����s_<|Њ�F��;��r^��kȊ�'�rU���T8��v�gnFR�UT
O�� `g��.������]���z�������Q�s2��|�q�c��n"�G]��7��8�ȟL�Y�t��ov�<%2��rد�sp'bO��c
>~�.m�z��[5ܷ�ª�Yg�>u&l"x�Ľ{n1'�/�,�,�e[�NJ����O������R���^{�匍��
�F��F��޲�_�~�����@�y���cbf>��R�����q)�i���W�֨�NAz3V]��E��4��`YD^�ƚ�57X�u�յNY�Zl��7@�8�l|V���B���!_Eإ����"�\�iq�	�?Z���9�#ӡ���9y����IrF��z�l#	#���棋E�俔ʅ8��Ƌ5?�Wf�G�?t�L��2��nb����*">��a� �\���< V����f۟�@h��I[��(�J�ƺd�(Gj��B�_��v�K����B�����b�L�ɕ���5]��G��4�	����p{'lק�Z�e�9����?_L��Z�$��hʠa-��9�.�qH�.�����3����&�L�hkp�Ԋ~��V���Wq��Ftv�0o��J�`nw'
˯*��	<
h{2�0bE�v2��]j�I��i���!��V�����<�`�_��*̾�ț1��MU�J���]��=J6V`m�����'u����S��Z�����jEP0�`p՝�]W�������h�!:��5Pxz`�޼&>�'��"�Z:E����\T�:��J����i�Ma]λX����>�}q�� Q.+�H@S�ɕL���:�^�#�4�e�.+��s�h|�'T叞�����AJS��x�2�p���?7fE��zO�=y@t��}����ʘ]kY](\L˜��轰���&u�ُ�);��"���'�"����Z�`��}-11��2�42GJԟ6F�U��䫮�4Y*�H���ز� ��
��޽{�F8G�Âߎ���`�)��ʻ	��=��\�'_2��t����ܫ}6s��!��_d�|&�� >}��>���������7o���f�S�Y��<�x���cP���Qy�
���%���Z��b�X�6����d�����/XP◇룇N��s�	r��aWu{ۧ��~�@��v#+vO[ּ��W����9��vi�a0o���@#�qwg�B���!��Q:����(G#�Xd\�1;�z�su�xI�f��D��d>a�Vv�|ɦ����k3d4��u�P��CP�.��幰�Fj"��)�u+
�����cGC��ݶt�|�u���*V[@~�A9�2��%_#AG���GkQ��>�TZ�t��dU��6�}����1fhOӎ1�O�V�ˬ�� Z�+ތ�J�`"_�R�S�뉊��qT�
�P�%A�5�\#a�ʰ���$�)��Ƽ˔����
w`��M��
�{�\�SǁG���#�j�*�,������F��$	<l��ͽ�s�7zޕ��T���w��]fT�e"��S��Z%��Y�P,�m+�RSr�#�/�B�}��Cg�S�,�(Z��x��ռss\�l�>���]]Bv��l9>�y�ih��m\��V
1����'��~h �/�2�DSD�{|#��9#�r�u�uS"COeDF
��dJ�m��a�9N{��}Wȣ�����j=N��.����i���\yۈ+M��W����6l^��]�/;���+܆�r�0�~�}���v�|�(�RD=8fk)���u�>���,�%����@[7wO�l�e�vJ���Ƭ��#떲��0���j�Q��d�~i��!��hy~tk��g/�!��FD�����=:y+
�G���pmI���/C�ћ%_*�U�.��J�
ӆ������ҩq�fŽh猾���U.��>��B~xG��o�����d�F��PJ�r����NX�������^g0�s)�A��;zr�6!!��y��qfP~.�����2���\=����D�h���Vҟ"���3��5�D�'_��ؐ�w�8�Ԇ�>� /�~��~����ҿB|�H�%��!Ӏ��I�����B襐_���D�& $�M�R2�XK!4[������*�ik9�`�T�#ay��)�=y\T� )N�W�+�@��~C�����6��h��Y<>+����`��V��nsrQ�#��oy�3�M����ycұЖ1�%�B�7�]�2GCP�-0��F'`"��̼����-��Tw#^��f�ա�G��R �ظ=F�&ЋU�@r�׉H��L.�~>�;�1�����\��m�c)
��A�L���}	ۤ]d��S���H�D��^E��+���^NJ�M�7�4MT��R���F��/���(����J�O�q�j��;��/c�R����nxH�i���� (�T��5q��p�t�	��E^};��)}�a|�~��"�F��$�vF
8�C!Z�	�rfc���h�2��l�`��z�i�u��T��fI\�pc�&��o,cI�ag�.�)�(���Q|�!Č�刷΄z�:�U�!e�E�	��wK��6c7�Y�͵� ڽ�!h��Aq6�����Dªa��ɘ�͖�bůU==�:�O����THV= *HV�f춫����؃��bk	���b�j��X}��<$��&9�D)S����W�̙ݳw��'��X�D���`���;I��̄QV�mn�AX	z�����κ�FӔ�᤾X�����@1���_�����tؓ\�2�p|��pHһ�;t>���<E��~�^�A��Pno����c��^��E��G~
�il~�A�R6���e���5�^����x7h�'3��h�����Q��Cׯ�S��E�vZ��N���5��^Gb��]z�xL"=,��	��l(��6�}.����!ǟ>������2ׁ�\&��r��r�p6JuK�.�/!T��.����~k�h����t��
V��[Ϟ����l6�zM��ʽЙn9N�l.��{e�罻OU.��غC�:�WG���]�8�������J~����� lW���"��g�T9H�G(􇘳Sh��E?�j�'�O��YPW�/7+u��N�l�n�s�/s��d�����M���?�O\�����b�aK�^=�v��s��Źø���)�y�����^��S���lun|��=���c�<����;�]q��<���A����<Z�
��qs��0�9V��Y�%�<�S�,J���tN�$+%�J��b�,�}-mG=Nʳ!�L�_�?@�䘜8�c8M=n]��B�w�)O�E���wւ�d��G֠�W,��ܽKw[yrb��c|	;HقZe���
#[�d�hQg�QP�F��Q�T&�7�9�6��Wdg�����xOӘ�l����q�]�Ѯ�V�����Yv>��F-�]e�x�*�!D|��yE���>�X��T1q`%'����
���D�<F�4J�|�~��H�z��l�u~N#�O J�{�"pW��'��"sF��s����	,�����3ceu��͒ȴ>Iz����T�_7���un��GP�����e���Bj�h��x�#��Dn:��0�C�	?���C~�Wn]^էm*�!rB5;yJ0�b_7 �Z �h�9L��r5��.a��C����P`?��$p�u֏F����0��~@4�6ʬ�^�o�"N 7�R]�e����m(ZZ�]�!{�+���.)ٛ�E��&7Q���gX +��ՄK�Էkh�'���ҫ32RG�f@�ћ�6ڃ�8���l��ES�Dv�iE��-n�B�_b��$����m��&��$��8I1}R�	�{>K��*YΖ�Ť>�Dx��d1f}���!��
`,�X�'i&�1�"d?/��� mQ��w,�龹�g����v���D�%�<	q8J���WS����2}��%-o�ji������a%f		�:QC`����w����ѣQe:�kp�E�a͜%�v@����q�.u�ټtํ|��b:w����ݘ"g�Y��Yi�ȅ�p��O=�.&�a�����g��U�~+��*72Xb��cT?ry2�ֲZ��n7�/ߩ�Zv^��ۋfDa�7r�=�q�}���h^�aЕ��
[]kd� /u�����8t5Go���ɬ���?��uzI��yt�S֧N}r�ssG���f���p�`����伯x1���Y�kjMK��瓞��+ �f��Jt�O��rb֙�Q���^��;pWb-��v�1�N$un�KB����V���{�G�)��$~� �ub����J�F5�,J�TB�^VP�6y�~l�=��[h�u�IP�(�6��� �T*�����܄�S�l��hЬ�������������Z���0,l��K��c%C+��u�w^ݗ���rerL������&�W��S�=U��O�1���/�}�<�2�w��²p��z��l4*%*[ք4ubl��djH��h��Tp�Y3�w^���i���M>vG%a؎}�rK�����cq�K)����9�]�.��$����h'�~���)�ƕ8y�Qu5x�u�(���It*]Gmo,�����_�i�yBV+�:�꬐��C���{灗�D�Qn��y>���h�]�o9�d O�YzE"Ԋ�J�{l���#��%>������e��!��>A�Y!�"�ק0��^����ubF�0��e�JE8�,7�_ޭ�K��h�Å�i{;n3�Y~2J��a�_���?�f�E���:2�v�����:?w��X��d4�w����g���T�u.6vl:V��\�.��������^�̪h���t�[0�!7V�4����7�\{*��FŖ��M��j��Xa�\�l聯��s12��p$Y�?v7��_bF���v+W��*y�������ۅ���iɬC�!�]��aVdJ�j:�L0Q��Ҳz8Z�9z^���M��(��Lb����5g��\��΄��BT/�_��Ш깬�4��Y�d��T�X�̔��p�nBs+�	��4���&QQtPZ��c��I;/�`^��N��y%�q��0h̸M������aDR��y�h�S'i�/py������f	�b?z�~n�FB�����N���?&?D�;��bCf3sQ{�'Q+S.��v�<�
/��fb��~y�E�H'���L&4���Fq�/�k�P��(:���G�z�{~��4�`*�%)�����"#��q;�^�&�����:�mljM��Yf�����4�{�rv���qX��T�o����ki�.p�u/�&�&Ԗ����i'���_T�-�ȳLr���w
�s�ż2�v	��i�ų��,7)��+�T@$R�v�"�Mp��c�Rcņ4U��"/7�f�����D�Z\�	'ٌ%5|0���\�y��ob� {!L\L]M�L��n���6i�-t�����<�ߓ�Xa��4.
�Ѻ�C����.��x�e��E#���e���pm�
�r�}1�G��C�ҝ��0ֻ����8���-ki�f,�֡9x�ԥǟ,�+�u���A�B��B}�$�Ȓ��0��AEF�ʊl���Ze]�Lb��8B��8ݻр���� P��D�eu���@Be7hQ�$�s�xgJ;���Ņ������/��_T��l���ބ_0�P@`�Zm�O��]D�7vb��N���=6��Լȼ6�p�kV�\��8Tw'r��s�p��K�vQ��	ri\e��x�=Z�2�V���o�@MK}�_Ѝ�� E��M �� ��מyk]��K�>�SLv���:,�SGn؆ǈs��R�dG^`J��W�!���U��^�q���}���D&[H�;�h��&}0�w�SJ�/87�U����S�_6ϲ��X�8Ac�>��Nre���jX}�cIO}��n�ȹ���Ă;З�j7�$Րu�|;�� ���"��j��=�V���%��X�P"!-�;���>��Р���QXڏ�;_��R�̒C)���0�����`2LJ<Ro=�I>9$|jYư��,��D�p�[ 3��i;d��+b��˟���.��ѧ����lm0��RT�Q	r��~�*nu�p�Y�s.�N3N�V��u�o��P�2�c��+�og��2R^��
���5�i�&u�de�=��c���o2����<C��ĩ�"��:wK�؀�& �z�yji��@�KF� �s,��U:Zk�?�{B������:��q�7���}C�v�獖g�䍩��O�J	��gLܡ+ O#���Nu����	��O?Gw�rp�	��,^�/nD�}�L��ͷ��}k���;�$|�>1EO�0���� �Y�ಂ>�.�t��j'�X�']�]�Wü�)�++���w"��ҧ���qd)p����S��>�;�~ð��@ү"����T�NM��YφV������,��ώ�Q�~��nզ�b��R �{��-�Y�Y=�̶�*�%���h:7�k
�d�_?����D(٪�^S���_k���,$n�F��3W�z��6�,��pA��x/�s�W<Hf���*H�v��E�鋼���V
��Tn���搀�=W� <�Zv|t�}� �5�wjK-@dc"fNIZ-H��l��l��$��S���VT("�eo��n��ɽif��fo�F&na|����"F��y�D�l�<��k^X[�����#+Kj�M����gH�D�ht�(7�W�v���4�M,�a#�����jIk��A;;�i!�Ÿ��cr�AW{8���Y]a���j�����п�����2���ѡ���J�3�)�rڇGG��J#ֱ Xv������d���=�ޜ�������{{�����l���d���hȲ��`�Lg���a��qg�������6����Z�q��/��pW9I�����[f{�p\��01�|
�n'2�\��~ڱA���-�<���<r����^*[w�4H\�Z>#�2��t���u����&ӆ��]^����5g�����2d�_���nKA0_+�����]z�-]l0�(���m��'�湱�� %��"&&}t�^�Ǿm��^�9���	N΁y�}aO`17V�pak�^_�X$%i�m�f>FK��΢���v�Jկ4���g��- ���9��t<Q��KCzv
0Z���ԋrt� %�:�e�����Kf��
��Xu�tj= ,�ф�7$��J�߼iu��S�]�4�oVT�(�x�P�i|��|�����L�[2[&�r�,���k!���FQ�ʶ��V���d���Vjճ�Z2���/���A��P� u8�G��T�vDIb��-7�e|�>���/=���Ӕ����G���av4(������q�呛�[�{�+j���?L�	
��.B2�����l��zyO��vNY�3���L�����t�w�~XT7�7�����.GR�~@�$��:�'��"�,ζ�e7��gp��0�e)��Ssq�V�&�v��f}������K��;�!�� 3���{�����#s#M2�ý���`�B�k��0Gd�
�A�CȭN��m+���B�!q)��7ڭF�����,�3>�����"
;# f������^�沙u��Ü���܅�QU�&D�]�
��ЮJk(vpW��#�����\��h��ן"��l�N^z��=���c��Ѱ�=CJ�;�|���ٞw�YS��{ ��/���8�@;O�S�@Hl�R�w�j���_/0�|ح��"Y�=���_��a�)T-]��:c�X׵gSR�tp}��Ӣ#�u�X�.*~K�N7�������Mgb���ό��?�rZ�c���Lv�}�%��1������E� �&AD�U�c=(��~k��گdeP!��	��b*Cء�@ ��J�k�������33YPh�W�!��d��#�T��j�H ,������0����-lP v��5mu�����N켳�L�E0o��K�?C�HK�܁�
6��B�h�/!u�f��D/�{���@���Ph��h��I��ݨߛ�{N���AX��ԼS�C�d���?���L�,rg3vhn C�~�]d���d�
VdY YK4\��vgo`��%�D���H4��;�Os ��bY%�	�z~���0d���,���P�h�W���h�Oª ƈ>���&/(����� ���]�h�6�����@a)ׇ�]�U,ǹ Os�L����빞�bPHE���-�Ep����-S]��e�E���Ή�݈�:�t��0?�o�����*C ��Sx��G�ࣟ&֡��������ȏ`����c�x�A��>nS��F
�C���w|�Dۃ�7�_�����hm�U5�dL�M����+�VɆ��&�)���db*�d��no�W}c��)�|���# ��>p�yu�q�V��"�"�H�$�B��b@�p"�O�,�Ϋ>�%&(���e,"xL�QM�����a�;�����u2s�Ř�s�G�9�\�I[e}��&L���-Ͻ!�7k�4�R�b�:6�<Z�`@��Ku�N�B(�)����l_#�;U��|/��'�y�*?�6���j�:EE�epu�d�gԴ�ߴ��wmls�YĽ��@W=�@*s��s��qc�6�1̫��d��gZ�X��0N���=�����΃W�z�v3/�oi�8���|�l �.4�R��&��CW�݌��*�NΤ���,�m����0�����b���%�k��2�7�����Dhc���[��ua�/�f�&���y4T0����d2�RS����� g>� ���t@�U�Y�(���$=_�k�ػڻ����V"բ�B���(�B���9���K,��@� H�mo�=J��H�9*</hQ؏@��y�&vis���rwO�����X� b��A���uCdN%��?��s�t����J3��0Oo�@MpQ�ɺC��%'0�Vm҄z�(���z����	�F�ẈHgK5����}R�q�y��b���7�[��g2�b����j^����6	1���0TN�\[S�D*X����л��<�6�2�̗�C��x�Xr"�g)oC�0=�|0����q�S�j��%���s����ɮ��p�ō��q��J��.�3!nR�F���CO�����(�#�*�1*��=���R�ޘD���L�R*8���\�3!�PY�M'�pʤ��X<�H$�����4P=a\Ʀ8�N�{y�� 3�u�k�����@���WE���W����|��?���]y�ېc������!d��-Rg|7���@	=C���I��\��)<N�6 n,;�L�n{Lښ	��s��(j3F����$$n��S.t�{c#���2�C��P{F����H��IO������F��W~S�\,m�����TE�t�F^���,��m�g�X\��',bQ�{��*I\�r���R�3�d�bPB('�jv�ʳ�#e�qV+���;$�s	A귡���V:M����ŉI�Ȍo3���p,�Q�_��i�?���3��6J���-��� "4)����<��$�d�����9�P�@ȑw��S���C���l�@)#�s|��ٚ�*:9�* |l����h�jb��ȕ�a�����GQ���R)��v��s��#��ɬ�c�1M�ɓʷ�2�$9	 ��#�QWj�Ȗ[p��1������?��L�I;l4��}H�n��x�2Uغ5P`���������m�Oo;�o��b�;���<�ț�;g��� ���r�ۛ�_�u��q����.��kпS3޸� �$�ܪA/P<Q�<`������h�101V�9}��#�+�{Gw����?3���;�HI�E}�� ��,�w�.^���M�]h$���(��0��Mi���O���>�!W@+pC1��ncn2�Q�0�*lc��+�u����m)}��g`-��a͊*:I,p�0(!\�J�����qA�ҺE�wM-�����ׯ���]�}��z�֓"̑� �B�~}L+��<���VH��ܭ?���ВjL� o����Rt�C�3KP6�0����A;V���0��dx��u}k��9�E�.
�Cǒ�Fe.0���!�i��Â� �;P�5$x����r�sq�~T�c��G����������!E�*:v-�tR;�\,>�}VF-�Zυ7�0�SR<9���ժr�v(�-�3/����8F��4_��C�q1��͜���X�Ix��6i��.X]��Ǉp���L�3�ؕ���$�o� 'HB��������-���K�J�����D
�������Q�W3��5a0`��ޙ�5R����f�����n��D��9O�r);G����RF�c�xx(�/��j�Q�Wm{*�tcäRD�p��^�9j��ie�ʰw×���Ԯ�CJ�&���z�~�g�͎o�����vA��C��3�:�&Q8��V��avTI&�ff���'�,ێ�2wi����,S%+aH	d�Ic^ˈ�pă�No�5aҨ��؄o�b���W�昁�ȼ�k���j$��b�^��d�9V�
~��/h��͹�T�1}�}�]����Ծ;���"s1'��	�bgN�,�TAﳆ�J�>}�.�:��]-"�.¤�,jtv�{�:P��Ol��,��T5k���I�g8!0����ŸD}��4 ��>iQL�6���6Z��M��/�`�o����X Z�a����Oa�܅ /f�[��;�sL����� �D��uo���S�F^;;C9�6��jf���о���&���$=�n�T�>U3�q�SoMA$H#�6����H�h�3p�Y�y41�E���):趕/��7����h��$��R�h<�?N8ϴ�&����Au�N)�EX��+=`�7�W��ڰ}X.��Kx�Y�q!?��9Y��ghx�!1�3�@ÎJ6��I y�J����S�O���%6m��d6����q2Ñ�)�	@�u�ÚV�ND2�d���E]o�dl�v�.��ZQm��L0I�܏PT�aZ*�N֣]D`(���pߚ:�DR�t �ȕ�Az9�H��,y��'�b�����$m`�4��
镻7[���D�i`�H+(�&�ܝr,��ʔg�����Q=J�6!m�F�E�"�� ����/���O�F�¬;��IiF��x�6��7���x	�ȭ�%��b�W�|Ap �.�|��#��;��dAq�z�z�����K�$�V0��zv���W�J%{ʷ	���ԥIl��������5o�m��x��\��Z���i5�|`�͢0wђ=�"��ю�!i-qS��e���V0|],F[���P�A�Չ٪g�3Q?�M1���L���`�U���������*�����6�)�&�${�������{@�젙(�I�����Vn����І����Uu�O���?N�<ե����a����cq#d�ҍ��
����LJod�d�M�sn�; �ȅ
oO�n3i�᚟;v�p�
��!�3�q���c�;u��]��èԀ1�8A��5}hjýR {�z_�<��+���5 �m|�fs��z��F�`3�A?�p�]�p'�By~X���P����e���i�Ĉ�Q��]y�LGʱbDK����O�6����g.�'AP��~�x l��6 ���w��h���4���Z��bD�56e��lZ����"��|Ĕg⇥��LN�ɮ����*�"4(@�̫v�����oZFI-�잼��Z���~�ܱ�nG:���k�DE��0�jt��9稏N[��m-q1ל������/g�M/���j�ߌ�����l�Jaё�8�cL ���"jk�^)���lp"�l���쨢w�lL�v���ʥ:E�ߩN�D�$�#�5��[#GvU�?���pJ
�U�`�pɞ��q_�

tC����|�	�J!um;Zd	����w���@Qs�M�E�/��(~#Ιڡr���q�ݡ]�6ϱtU�	�IFbDo���U�`U�~֌� �,���_)s�݇A�
�Qll 9��`�1��]n>��qFb?ߡ�B�9vRzumm�_	��U_f'Y�ix6Z��t��U��?�����;���4szC�[s�;��ꌗ6��2pve����U�Sd3N��.=��F60��ˢ�c7\��0����$�z-Wӌ�<����-ő(a���?���j�/��I�`&Ζ���L:��/Ami法�D��������b�O� _�][S��)�{�Ĉ���"�1���*�Ep�(�L�vR �86K��Xτ7�I�d�S]�n��+���ø�W��P-b}&&�}����#��-<�R��
	��>��2�%� ���r�/c���w��IiT����wP(䎬�US��0�b�	���J#Z���¹��*SX���f_�5t�����(q gZ��ʢ�j��)9z�b�C�������ex��S���r�� �YF�o�+�{��L�z���3��t����6?��u�2m��\*EB&Dμ>0��R9lQ�(�?���ߺ��h&���H�0�K��/�_t8�v��s=��ɔ@�k������m]f�L�����Pw��XB����v�'y�!�/�-I��xEZ
�������0c��E��H�G�.�)�*�a��f\v�g4��
Qﳬ݊["v��vq.8�6���[��������'���� z��M`�t���1���?��W�RĞfG7�f���Opƨ���v�$Pug^�K���� ���\$�+$6�sO6?�̛e������6��;x�I l��hã����/Y�q�|2 A�`>�&����{���1��2�R�v�i����@g�I���ǚfJ�G������%I�ힻr<	����˳�F�ˈ�6$���'%v�,>`G�Q����bLd��SB�As��?�l��^��n�!M�'�u���3�u(�0�C�l���_>Y�a璋�L'g)E�)�AS"�'8�Qab&ki\"�:�_S�H���j���B��*��;�Qa+:vk�hL���Ϣ���+[V|�r4-E!&��~]A�v��aGd	%��}dL5J=�<ugN���rؼ��k �*$A)I{�@��<ZCck��Y��R	<��h��o��T*8���(]֞vv:�L�_j�\f�k氅�k�����#�z�ep£eܹ�\ � r�I���U!#u�\R#9X��xsd5vq��41��JnQ��<�'�i8�m!恅�6��qr�GF�]��3���O�����,��F��;w׵��R�^V����&�b��ߥςN�˙�S�%D�w����#H��@T�a0�R�tH`�yR�;�J[�������?�źa�A�hx:�'p[NÎA�c���Ǉ÷��+�Uͽ���$	P�Ip\̍�F�9�p������	ҽ���EVap�H�Y���/�s�׎��]�R��9��G�r���	8�7tU��7�C���kP`w��_�4>�A�׊ 
�������kH����y[������*��s|�57�@�KX%��`���r��a-tMl����}��]W-̌65C�P���Y�8h~@��+�G������B
����2˷|@�=y��� ��W_�v��jӌ9YԴ����Խ�E��o���'��6���%�xs�r�W�w�	���?�4^+����}GB|���JuȢ�4I8�zစ��(��Ղ��.��0Ɉڶ��fq���V��M��B���0D��%���y��?U�DK��9:�hO�~i.��;L�k�2�w� �kӌ��m^��.������b�<�eM�g�l�}x��@�*��Mq��l�u���"��=20�YKưt
�@�xd-v��a�xdr�.!A<����K8�I0���r���*b�N �	��$_��-<�`ᕇ��?�)�8�x�}�R�Q��Dܩx�{�Uv�泂f���|Nj�r�G�bK�Mˮ	IC2�vS����׋"�` 	���=� �2��/�L6�>�J�_�2�������%f'u΀y%��ۭ��Ϣ�-���F�z�#�0�
��K㞥�ք�5��zd��`ېCڜ���Q+�
��զZp���G@T�"� B��q�z���<��`���(������t�����"��.�N@	��+P���0z�]�QK� `�p.nGŵ�y�Ogk![�������Yh�Ѿ��Ec�	�����6HIO�x�h�Y��HY*��/��%��$�ڼ��A=�^]��F���k�p�ɚ`�� w9��uPuU{UJtp@w~���22�+�p'َ^aWĨѮ��3��e���*ů�X�7�%IQ�d��P��7��o�B�"�����p�q��Ǝo1����O,Îm'��<�>�v���(���(>�ͩ5���gc
rʸtx��ׄ���,PѶ��+?�jdQ���e)c� �J�U��J���.ͳ���PG���p3�ߎfw��2�>���X����������}��oI}�8i�J����<J�=�IyUB��=~�ً�U��	�GL)ǰ���QDp����x�E�=n��3�{�>�:^-�����0a���0K�A\� шTN�����}�pJ�CY��=Msٿ%���R����S5n+�5Y�\�o����]Oe05��� �跀=�Ȏ��S�Z��ŕ�};/�T�_%�f�Gûu��9�|��%�Բ&nH�qF��͕��*
��v��D�l�DR<�>P������o�]�"����~M��F��9zD� �T�tX�;��&��R�_�zG�r��i�jĘXs&|EWB�["��b��K)���k��Ձ%�*�¬���$Zd�'���YkG�����Jhl�8;�j.��/��i6�M�Ȳ���p���E٘G�[l�v��֝�B1g�x/0%TB@~©�9��k_m28��.3�Ι�\�`o�� ���ےRabC9i��(�Z7�.�=�\!�2�&�����E��4���ڔ�&P�h�J�yOB$��������~줁��3Ɩ�2�^�N@�����h�:ZF��.q�wL��wU���n�\��KDD|?!-���.���by�ɚ�Kg�D�|T��+�������K�C�C�1��H�|��so�M���ߴ�>���"X#p�F������X`~��n4�r��~A�w��-ZJd���Q���u3�X=pB_j?\*<<2��Dv$����ˡ���f�"�u��p6�v	&b�.P.b�cݥ6?�N��kMqI a0�
J���F�B{sO/"�ћ�Z��6uM�?��:VT��C���ޓ�MD�U�^�B����J�����9z_8�� �Q\VD	A�97\}M�s�5LwDj���Q���ZU6V����8��YЁڕV!H)VҎ�M)h��'y4Զ�8Mu�jI�;�O���4�1��P.w/#�C"W���Z���sY���-��7����N�=@Y�_�/u�(��yS��t����|��fO�X]��K�od2�.�H���d�X�'����SQi�����Ilp;=p�-������z#h�,D)WK*��KY(U�	��6]Xh�����d���c�@g+�?`|&�u�TO�o���q���0Q�8q-	PX� �
�	M�A�G.B�QUˍJ�����4�����)Zʥ�������TA�S�77UP�՟�;�};T��%��#������@��~h�^ԏ�&f�#a>@N�PN3T�0��:�dm�;e�M6c��r!�?���t��E����� DdT��u�zRv3��)U#�ZwU���m�?{ǣ�Br��/��Ο�����Z.BMࣛ��h�,I��G$�(v�j���G��*c���kSe�Yj�AB�*��^eO�H���� ��Z���3��h?��[��w�(ӥ��ä���s�3T:*�M�U��E1��0:�	�켸:z�lr��5�*�D�U����!CU�]\J�0F%|��6�$`�W�a���2���#���d�ЙG��~P�7��׽U�)��g/��f4C�W���z gV�m�
K��a������8�-%���Y���q����{<	J���َ�Ϙ�r�5���t�
b����&b���u���dJ|��l�0��$@z��l�r-_��i�����xj�-��.�t���L Ff� 0�<po�<>�:����K���M�/���1#In�Z�ȉ�T��k$��6$FЍƉ-�dw���1]��B<��L�/�29�cOo�Ⱥ5x�3mL��2��F��](��v�����j��xc��xwc䰃	�
����\G˧
@�[�Ƴ�j���ߡ��l���x�l�����_������iAQ'Ȉ~'�]VD� %�遀�k���Б[Ƥ��u+����2����D� ��&��aԉ�=Ӈ�x8%Q��y�+��G7%H�6#* �|���bfɅ����zU� ��Z�g�o���s��BL���~��I7]e`��Y�u�uVa�D��h#QC����Ź��6$f��D��~��~.������3�y�N��\��U�5��XFp=��=B�ޒ�zq].�YS�3�7���@�\�5L1�rd�;ct��h��GΓ{>z(O�K�5������*��%]�~<*HK�$(��\��⣥{7Ɠa�k��v��%'��=���d������9�}O+��F]����(6M{������ c��E!�,s���"��E�97���_Dcj�,��maㇿсiox���.!����2��a��]D��L	ޡN愵����W�q%<��҂�lpX��J��T#��i5�'�:�ov.艎CbI����Sͣ�|7�>�#�i���Q���Q���8n�^y���w�0�:rf!�n� iq�(�^n��]��|��F�m^H�����((IT;?=!<��A�����uӞ�=�"M�
ep�Bq�#��9h]&ܐB!T81o���q]�1A��[����J_�
���N9���s�e�ʒ�=�V?K��� E!8� 6�;��H0V���Gb{ȣC6R?ʅ讬�D�� ��?nt��ң~���o�� x&-�pT�h���M�N�rX�И���C+�N��>ڋζ_~�����4=9������m��Qi�vOA�ԕ ^�2��vQ6<�"�sf�w:���L�!�U�,������(�Ϋ/	@�r$J�E�$ړ��P����h=�	��x��t���a%oVcs�]K�B{f����-�p�ܐsc��~�ǻt*('^}*�h��B���X�7���4��SݛJ2k\�gzV7����ڛV	��uz�h��P:@H�J��'w���pM�	�#�7��?�_}hK�I�=���ړL��5��G=��O�xםe߳ڧ�l�Ӣ,�x�j����тZ,9�'3�H� Ǉj5}��YJ��2b�+P�����h<�B䡭��ߡ����Z��ژ��}�l��\�_h%04���o�y� Y��ާ�X!,3��J:�ǁo�ˑ&�S	��<��d�5z<<��!k�m�9�OSa�C����<������g5��y�
@ nϘc"�L{������Pԑ^E��p)�CF[LH3����銀hI�� '���yp┿��3v�z�;�����Mwt���W98�a2yC�F�Ƃ;O��OQ]��c������isԀm�VJt]�Uq��������j���s�/L��5"n5m7tT��da%I@���G?so���� ��:�c�Jh~���3�t�$��_#�0rG��$����g܍����XU��F��V�5��;~�1�}W1�@��87Y�Q�_��J@�OKv�`RM���(Di{N�g���?s�l|[qخ�����I���b������cBH��|H�����6�J�,�n`h���)���h>�ˌ��{}*K5�_�s�����G
U�83�W8���
� ��`鳼�c��$g �"��O)�M7w��nKa���7�m�gmSۖ.�\�D+r�ߣ�٠KQ�W��GC�!�!s�v@���	ՒS���F�P�+���MX(n�:g"�||�+YZ�I��)��nB}��^D�$�.��Au��O�ŧ	�	���z�|�@�#�*�Xw���Y��b�i�'�\]�5���V�D�![�\�����9{9j-���qe�K�(b�*���@�efvb��͌�����,n}�����Z[�e������ǞF+_<�� '" � �p��T�I���IeL���
͐�1x�9�u�bΥ�Q�Dg�h��5lC�2�
,��lc�d �,�C�ʞ�&