��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.�ܫ)�/ ��rbm	P���ע��j$aQe��d�����![�1�Q���&GLM(��;$���^X��H�U���-�18;�ޑ�Q�ahABA���M��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�F!�L�� �ٵ�˔Ɖ��� D�[\��:z�^}���8.j1�dLT8ͧ��t�%��P�B�т�R��U����-|�8�3�ԣځe'V'ޑ��s2+6`���j)L&��؛���kw���B��(�2r� ��֩�5
�~N�۱��]�tCB�rZ�4z�5��o�Κ�{����?��>�4WyD#;m���Fh/Q���}��O�aW��ޒ���
�E��vtb���45Z�2����;�9A���}�����I�v���[�
�<��H$9	���5+��I�����u݉Ll�c}��Hf�ѻ{�I��3N��bd����k�F;�E�\S����Ýi�I�p���Q�]-���|���3*
����D�d�D�����k�\ ���#�kX�XV��pBY��c������#� ��+C�Q��� �<����c��<0bIx�<3\�쀋��.�-\g�
��J��L���b尨q�������*���s�5#��э��$��C=֌S�2'��6t��X+F+��o�pQR8fp��w��&Bd�o�CZ�!!� ���M[pI���W���z���o�e���;U�ҙ"I�$��z��GB��U�k���YʯGD-0c�Ed��}i����B����H4O�{�U�m�9�P�ΣR��S���������i`�t��*7�/�2̑� {��nZ�e�1&�G6�Nd��2b�g�R4 -B~�t|�De ;q +�U�����C�Z���[{G�(��"E�d�ݱ�����\�n��w�k1�k��20�t0�Iz%졐ϔ���Y�3ub��U~����3�d�oB �n׭z>����k��^h]G��Y='���(�m�/��)�6Z�e~�R�(GJ�;�r�U��Z-=}R�����9�%i�Ǎ$�I��m�Y���]���j�j�
ŇO���Kf[O����&�bO��O,�>��;�Kj�#��	?خY�%�T���C(g�)�s��d�����`�&w����,�{?ˠ7��i���ף9���4��Ard��'Vp\�G�����I����v�)bn��nc���� ����(j=r��п�͘�$)�|x��Ӟ���C��4�Z�跟��uPq�M?@uǿ�z�N����c�:#">��ɒ�d��znU��w�<�`���ߙ,g�>
�k�Ѕ,�"�w_?8ݠ`������L���텻T%cᧇ��A;�X�˕X;�J)����P#��i�$�v�~
Q҉���ȡ-�.اdQնg�9=�Q�Jy�AɧS��PA�H������q!����z��[��<�4w�vs?<�Z|W͛@�� �g���gP�$в0��	mOrl��%9b���B�Z�[����f*s���d��Y'f�[�5ܸs������5'4��g����������WP[�i:��6GN�4mSť���XS��� G]8<��X�+�O/�����{��\1�s���PPW��5G��2b�ys(���I��l�	��V�o�]>q-j�������4�t"���<0����Lj�~W��ɀ|����9�j���h,�g�TDӻ�V��,T�� ����~�Aֺ���5����XtC��D=��2�HH�i���ALS���V4�a,�h`6Q�#2=x>k�~����B�a�,�z^��z�$�3p7�:UӴ�ЙU�`������m4x=�/4,i@E�}�(fQ��JF0�z
ȳ�3C+�㶰=]- U֦�(_;�±!H���by�
�c�qB0���AM��r,�����
X���c�M���m�OsR��S�h{����T}�7'[#p��`�"W�����+X�U;E��	,U��#d{��9�}3>�ہ���t���0�be��y�1�V�Ƴ�.����X��L�i��B�(�� � ����qd�M�Ȝ{��g� 4U�	�ʩ�B".^���[�1�"�΃f���������OS�7o��M���<���]2!wn�K���˨�\��(�we�2χ��X���ջ���֯0O\�*���ԋ�E����x�����/��:t�h+7�;/��qNG>�C�@I6W{��Val%���=�(('��kɦ&_�o	T3�֍~���������s��*���v��޶OMUB�����TK������dA��v��&�ixˉX;�-�*�V����E�q2<UtX%����	��l�h��z�Rsm��Ƀ��C_���Bb�����[�
�r*�f^!A�������p���wXEՕ�b����^}����Y�j�F/�/�/s�2
�����;�Ҭ��]{��������$9L��Nb|�^���ֹW^�Ȯ��Y9`�$y�@2��n�����q�S��>��LjH�F���|����������|�oR�����8�!!E6���������ѸD�����7~��1����Y��n�6ʴh�y�ap�b�$�"}ԋ���zͩ� �(yԧr	�MG�.LC�*l���쪭�~똢���2����Q����
�°c%B��%��������e��Ir��A�.�N���R�wZ�Z㐌å�����ʍ��W�#ӊ�Ou���}#�
��^!�Җ�Mj�F�Cr(>/VS]I��_�o��X�	6� �S�$p��HV��C�����6�~sK[M��Acݶ\�xE?Ѝy���
�lΚ2�S)�ԽB�Fʋ����B��+4g���d)T��d����QI7���	Ѩ�X�rsǈ��x8H}��y�c��_h��N99�)�\٨�x�!,/3f>��Z�
A���R�i�ڿb�5g�i���f%W��jGY?~2�ax���!��X�iЂ"�*]�S_���C't�c�������^wvP�*�e�����}�CWb�n(����\�����a�ﮏk#vӄ5IE�9��B4cj���9�Qg��ٹ�窌�l�bN �(]��M>�D`�"o�2 n��ͧ�n~/������1~�D�QBՖp��M����T�T��E�B��o��"�t(�`΄�>)���½��kz��'[��>�B��+��U��>�[�K�Ya¡#⬰{
@y�@2�s�*�VH{��;u����G��z����F�SV9gл�[�X��r"L|�u��ǜ����/XiLQTͮ�2Һo��[ro�["����'ʾ`�T���Tw�CwN��t#uG�$k{�D|6�KJ�i���i�