��/  "�	g�Jp��kV�e��B��)}-QLoY�����a�fܢHVn4��wÊ���0�F�ނ�3���.��aT(�,o���|�����em���./�����.��Ւ�!��� �廉�%��g�]�Z�Zf�s�~�� �����e� ip}�mR���'I}�7P�:I�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���w7F&3<�*/��컆9�AGW�?��J����02�,�����W��ž��<�U�7��eJ��vWz�;`�¹E���y���Zj&��j��Ԋr�ߍ�l;ZU+���*g�I��D����SC�q�XP#�~�#���@w#D���0��u�w-ett�$:he��}�r|{����qb�p~s����7F2�d����##&���p��laz0Ą����&���3[�:�D��g��ΒC�m�����9���(E�<�7��T\۾�~���bC��>^��k\1����>s04�dx&�mf6����(�򃝩�U_��;�ӵ4T4��֤߅+�*��i��P��]��$�N�
xK�kޞ�B\)���O �ț9�]�'���$B?�>�.7���>��B��S��1�
���t"��:CI��\*��3�3ŝ>D����*X�L�U�&m�)�R!��+*z�Q�A>�����٠��Q�αV��9�>��`�Xԟ6�A�L�������>�e��n���(ob_�z�����a�s��E	������خ4x5�����M"�9���N5go�4�V���h^���kV��<W��ݽ���u�	wn,�D&����?�R��2����=U�3��YV%�犾淏+��ˁ6��#�O��&eP/e���9+/~�	[�C7R�-�C�E$�����Z_W9��M�G���}�"�����A/=�{���I��)Q ƻ�@�@�:*�*����ϛQQ���ݾ��U�VJ� ��`ܴp�?S�v���V'�I�^CJ$9�WA���|���[ ��X�H�\$�x�$����}> `�X�2��r�6��Ω�(��`_w�g�C�����|>�^��ˬ��k���&�M߼ӯq�>s@��;���cO�(0�i{��c-,*q�.$�0i2���O�(��t�,-�q=&.{�]��H|b�&J����3�
V���9��)_d�b鎾��"�pO*)����-�g��ƈmm��(��H��(i&l�>h���)�=b"J������ӝH�l��:���k����/���)�_�T}�V�v�5�)�����c=��(R�m��-��o�����$��wI%W��J/�$����\��$3�	�,d��a7�!t����&�T�������pw�{�LjfykH�y��o���Y�*<0yi�d�
07��wt�8�`sr�W/>ո�)�( ��FE�z�Datu6'�TDո+�V:s�}�Ϝ0��ҪY�ƻlۮ���*�A���Vcf\j�#~����|�#����o	�����c]�~R��7Qh�f��Ň�P��_\o�0��1AK~]�l~8r��b�'XT}�����4Er'�[#���g� �1�
����B�-��@�
�8E6�CO�Zf0Vd\÷���u\%k��%ᮛȀ�?U��ݹ�u�����;.�5����E��mK�̒;@�_!1*p/�¶�Fv(E� �q^��b�N�h��]��ͫ���_�O�&$�fk�I1�CCz��lܷ����K�HӗP��2�� �X/�Ц�K�by�H��u:e�'�m�a,|W騎N��ßw��� t��z^��� \$m��X�1�s��Gt$I~�/��2���T��=�� �NQ����既��l#�J�����1���Dv�R�����^tʒ�bb�Z�.��`>�A6� [�pM�>]���Ϸ�O�4�yIɍ��THy�)^�e����˜R�O���{��%��F�+X�a�wȶv���O�;��.qhS!.38�iG��1X��0�e�D��9�@"���sd����%2�
�ʦ5���:)^��S�A�B�ë�qLo]I�맳t�A��#$�xA�C1EC4�@|.���K�۳��h�4�fq��%LY��xʈ9	��m���2C�� �P'n@QB� s��ȓ̭�7�j��:�^���0o
(\n6eȕ5{�y�m�%$����ʷ_m��ű��E��{�%��%?^�s����.������G��
��y;ɡ&���X Eg�p'</�!��Sa�]�cZ\k��.�i��}ʋ�L +�VF���V4[>1��m��У}IvА����8��mQc�8���<G	�T

o��jr���p�,�x^� �Vn>W@�~`���������]N�	���Δ�u(f�4��À��k���@~\ -kM^��pk��PV�x���NlF��J*��j���C��<h��e?��z:�2��f��+�6�5�6� ������ٵ?�~4$�����B%
&^����KՑ��v��5|<Jr�n=NJf��?��Sdd$���bf[~��*�M,��W�;�UAD���&!/>��V���(��Y�Ja����oT8j�yL�j&�m9w���R���Wb"9�c��ɒ�)H��恏6�)��Y���Yy�|����/=g2;� ,jYo�׋�h�%�Ta!D��\�{4��),��1P�.�d(o����x<'1��-O2��4��N�ܹ|Kh��%=��Ǔ�a
�l�i��@��-+W˰YE�_h� ���6Q�~U��L��S�_
;hA���$�U�Byx��;��6]�zz�L�A0`�h]T�)����v�o���j<b�DϷn��Zw���0�.A��."�:OX��6C��:Tl�{XzL��ǌW�Y�&6�����������Ȇ�#��LS�I9�&hb�<��ȭ]A��&�ˌ�C{�4�X��]m�,�ʫ�fTh�c(�_����r�{�X���M�R�e�Io����//W��$���2�Ӯˣ���.IB	�K��XhY%����#�'+c�YM���׊�~p���EV8ZX����^�g���jIxӷy��XdG�����K,�+�k��֊���g�:���b����v���w�eg�@��F�`��A4�W��;��*��qCk���I'C_7߳2�v96(����hd�%�������<a8z�T$5�7��h����)p�Nҡ]��2���vp�Oڕ�G]�GՀ�Z�>S��K퟊Xv1ot��B������O��؁R��/�����v�>'%^��ln��g�vm�܂J���S�{�Us��d	"��㸃jx�����$.�9�����?��,�`Y��|&V?E����mMnK��˭T��4����Sf/Y�"d���T�Ö��喋h����!���U�D��J��!o�!�_A�n1,Q;�$��ح�픽���f='�$�� �?��"|���)6$�c2���Ooh�(fl�W�J�~<�1���T(ϙ���S�F�SPu�|��iĆM�8�:L���%�WШ̎;�d�ͱ���^&���/�'�Z@���y.o֬u!���N��E��nY-c�&���2GQ�Ow$I^�	�.q68e3"(ǚ��;�,rXQّ>��hc��7v�1Կ����ܰ��`�N���[[<���m��C��7a�����&���QJ��]u��BW�>�b=�mȔ�0'�Ilm�g|#-Dl�������bR��)��{ׄ�r�4�5�Z��p\H#�$��/�
@���q����=��ĕ'*���2-�-2�<���d_H5�<�����^O�t��2�/��W��h�M7�F�!��=�f9ļ.��_���9���7��E*T됄8�i��5��]�Rv�Ƣ8����e��o��j�k]�J������M�_�	��I �T^ֺ�O��SزX۪ZJ���(;��G�U��ϲ�	��ۦ��s�cs�Ҿ���}����<��F�侂ױ�
EӀ=[A*�x5󎓤r�'m��W����Z<I������&�Q��ǧ'qG�����Ts����wåQ��5���am\_ ]�X?��4B�N=�<�=yln]�H�̓C*���C��-I��g�:��y��ٯ����MFM,$��,�bN5�o,9\��ʹr�)/��_� `_	ʲ��\�P�D&d
��kB�?�Mw7cB�QÙ�)l��Pn}�}ڜ= ��'���A��-RSkJ��oE��!���W�#� ��@]�E8��d��A�A���PuLj�h�&h�mu���3;�;���/�I��{���B��zZ�wPȋ#� !��6yP���MbaE/��N�|S�h�`+�̬x�l<5�@A���\��i�at����?CDn����P���sxbι���]5q�����li����Hs�H��k�����F��~Q��C���V��L�e�b���ω�H�\0SD>�6�cI�j��:�R8��b��!��7��_#t����o��v%�Ә?,��)A���L>A#as�'�!�/��A���Y�1����!֋ާ��)C����aT�]&����s�v�|s���+R!/��jK��l�8r����@xx-�\2���쟖�3�,5�\Z��j�ϊD�bW�U{�����Q���בK�QF��%R�F�7v��3����,�a��vwDRwm���@��t�W��7Bw�g�)�ϝ���b��|�R�ᖜ�HZ
�)3ꁗ��-��+���v�����.�.����^V��GC�TJ'����\T`n���2�v�x��f���:ї�s�1E?P)�|g�]I��]A��[ӑ�wsCD�	�N)��y�z�+��X������RN^�����	���]�T1a�ڄu~�"�[4�Br�J��G�X*��JƄ?{���P̻3"�Ftܿ�����bܜ�jj5�0C�7K5w�<d�E@�؄�s"!v�5ɁX���`�*<K���P�`�7fl�d�n���P�+��|�E��Op&o�"�z�������+Kj�`[�g:����CQ�6��B,b�3�]w�b���I#�7������ϡ��B�ֺ�`��ˊ笑��aV�b�#>Vs�Ι;a0jn# �VZ�8��FuK�U���e���_�u���(爆��e���-G���^�"���5��`��-T�:���